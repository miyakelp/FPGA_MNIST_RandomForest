module mnist_rf (input wire [783:0] image, output wire [3:0] result);
  function [9:0] tree_0;
    input [783:0] pixel;

    reg node0_r;
    reg node0_l;
    reg node1_r;
    reg node1_l;
    reg node2_r;
    reg node2_l;
    reg node3_r;
    reg node3_l;
    reg node4_r;
    reg node4_l;
    reg node5_r;
    reg node5_l;
    reg node6_r;
    reg node6_l;
    reg node7_r;
    reg node7_l;
    reg node8_r;
    reg node8_l;
    reg node9_r;
    reg node9_l;
    reg node10;
    reg node11;
    reg node12_r;
    reg node12_l;
    reg node13;
    reg node14;
    reg node15_r;
    reg node15_l;
    reg node16_r;
    reg node16_l;
    reg node17;
    reg node18;
    reg node19_r;
    reg node19_l;
    reg node20;
    reg node21;
    reg node22_r;
    reg node22_l;
    reg node23_r;
    reg node23_l;
    reg node24_r;
    reg node24_l;
    reg node25;
    reg node26;
    reg node27_r;
    reg node27_l;
    reg node28;
    reg node29;
    reg node30_r;
    reg node30_l;
    reg node31_r;
    reg node31_l;
    reg node32;
    reg node33;
    reg node34_r;
    reg node34_l;
    reg node35;
    reg node36;
    reg node37_r;
    reg node37_l;
    reg node38_r;
    reg node38_l;
    reg node39_r;
    reg node39_l;
    reg node40_r;
    reg node40_l;
    reg node41;
    reg node42;
    reg node43_r;
    reg node43_l;
    reg node44;
    reg node45;
    reg node46_r;
    reg node46_l;
    reg node47_r;
    reg node47_l;
    reg node48;
    reg node49;
    reg node50_r;
    reg node50_l;
    reg node51;
    reg node52;
    reg node53_r;
    reg node53_l;
    reg node54_r;
    reg node54_l;
    reg node55_r;
    reg node55_l;
    reg node56;
    reg node57;
    reg node58_r;
    reg node58_l;
    reg node59;
    reg node60;
    reg node61_r;
    reg node61_l;
    reg node62_r;
    reg node62_l;
    reg node63;
    reg node64;
    reg node65_r;
    reg node65_l;
    reg node66;
    reg node67;
    reg node68_r;
    reg node68_l;
    reg node69_r;
    reg node69_l;
    reg node70_r;
    reg node70_l;
    reg node71_r;
    reg node71_l;
    reg node72_r;
    reg node72_l;
    reg node73;
    reg node74;
    reg node75_r;
    reg node75_l;
    reg node76;
    reg node77;
    reg node78_r;
    reg node78_l;
    reg node79_r;
    reg node79_l;
    reg node80;
    reg node81;
    reg node82_r;
    reg node82_l;
    reg node83;
    reg node84;
    reg node85_r;
    reg node85_l;
    reg node86_r;
    reg node86_l;
    reg node87_r;
    reg node87_l;
    reg node88;
    reg node89;
    reg node90;
    reg node91_r;
    reg node91_l;
    reg node92;
    reg node93_r;
    reg node93_l;
    reg node94;
    reg node95;
    reg node96_r;
    reg node96_l;
    reg node97_r;
    reg node97_l;
    reg node98_r;
    reg node98_l;
    reg node99_r;
    reg node99_l;
    reg node100;
    reg node101;
    reg node102_r;
    reg node102_l;
    reg node103;
    reg node104;
    reg node105_r;
    reg node105_l;
    reg node106_r;
    reg node106_l;
    reg node107;
    reg node108;
    reg node109;
    reg node110_r;
    reg node110_l;
    reg node111_r;
    reg node111_l;
    reg node112_r;
    reg node112_l;
    reg node113;
    reg node114;
    reg node115_r;
    reg node115_l;
    reg node116;
    reg node117;
    reg node118_r;
    reg node118_l;
    reg node119_r;
    reg node119_l;
    reg node120;
    reg node121;
    reg node122_r;
    reg node122_l;
    reg node123;
    reg node124;
    reg node125_r;
    reg node125_l;
    reg node126_r;
    reg node126_l;
    reg node127_r;
    reg node127_l;
    reg node128_r;
    reg node128_l;
    reg node129_r;
    reg node129_l;
    reg node130_r;
    reg node130_l;
    reg node131;
    reg node132;
    reg node133_r;
    reg node133_l;
    reg node134;
    reg node135;
    reg node136_r;
    reg node136_l;
    reg node137_r;
    reg node137_l;
    reg node138;
    reg node139;
    reg node140_r;
    reg node140_l;
    reg node141;
    reg node142;
    reg node143_r;
    reg node143_l;
    reg node144_r;
    reg node144_l;
    reg node145_r;
    reg node145_l;
    reg node146;
    reg node147;
    reg node148_r;
    reg node148_l;
    reg node149;
    reg node150;
    reg node151_r;
    reg node151_l;
    reg node152_r;
    reg node152_l;
    reg node153;
    reg node154;
    reg node155_r;
    reg node155_l;
    reg node156;
    reg node157;
    reg node158_r;
    reg node158_l;
    reg node159_r;
    reg node159_l;
    reg node160_r;
    reg node160_l;
    reg node161_r;
    reg node161_l;
    reg node162;
    reg node163;
    reg node164_r;
    reg node164_l;
    reg node165;
    reg node166;
    reg node167_r;
    reg node167_l;
    reg node168_r;
    reg node168_l;
    reg node169;
    reg node170;
    reg node171_r;
    reg node171_l;
    reg node172;
    reg node173;
    reg node174_r;
    reg node174_l;
    reg node175_r;
    reg node175_l;
    reg node176_r;
    reg node176_l;
    reg node177;
    reg node178;
    reg node179_r;
    reg node179_l;
    reg node180;
    reg node181;
    reg node182_r;
    reg node182_l;
    reg node183;
    reg node184_r;
    reg node184_l;
    reg node185;
    reg node186;
    reg node187_r;
    reg node187_l;
    reg node188_r;
    reg node188_l;
    reg node189_r;
    reg node189_l;
    reg node190_r;
    reg node190_l;
    reg node191_r;
    reg node191_l;
    reg node192;
    reg node193;
    reg node194_r;
    reg node194_l;
    reg node195;
    reg node196;
    reg node197_r;
    reg node197_l;
    reg node198_r;
    reg node198_l;
    reg node199;
    reg node200;
    reg node201_r;
    reg node201_l;
    reg node202;
    reg node203;
    reg node204_r;
    reg node204_l;
    reg node205_r;
    reg node205_l;
    reg node206_r;
    reg node206_l;
    reg node207;
    reg node208;
    reg node209_r;
    reg node209_l;
    reg node210;
    reg node211;
    reg node212_r;
    reg node212_l;
    reg node213_r;
    reg node213_l;
    reg node214;
    reg node215;
    reg node216_r;
    reg node216_l;
    reg node217;
    reg node218;
    reg node219_r;
    reg node219_l;
    reg node220_r;
    reg node220_l;
    reg node221_r;
    reg node221_l;
    reg node222_r;
    reg node222_l;
    reg node223;
    reg node224;
    reg node225_r;
    reg node225_l;
    reg node226;
    reg node227;
    reg node228_r;
    reg node228_l;
    reg node229;
    reg node230_r;
    reg node230_l;
    reg node231;
    reg node232;
    reg node233_r;
    reg node233_l;
    reg node234_r;
    reg node234_l;
    reg node235_r;
    reg node235_l;
    reg node236;
    reg node237;
    reg node238_r;
    reg node238_l;
    reg node239;
    reg node240;
    reg node241_r;
    reg node241_l;
    reg node242_r;
    reg node242_l;
    reg node243;
    reg node244;
    reg node245_r;
    reg node245_l;
    reg node246;
    reg node247;
    reg node248_r;
    reg node248_l;
    reg node249_r;
    reg node249_l;
    reg node250_r;
    reg node250_l;
    reg node251_r;
    reg node251_l;
    reg node252_r;
    reg node252_l;
    reg node253_r;
    reg node253_l;
    reg node254_r;
    reg node254_l;
    reg node255;
    reg node256;
    reg node257_r;
    reg node257_l;
    reg node258;
    reg node259;
    reg node260_r;
    reg node260_l;
    reg node261_r;
    reg node261_l;
    reg node262;
    reg node263;
    reg node264_r;
    reg node264_l;
    reg node265;
    reg node266;
    reg node267_r;
    reg node267_l;
    reg node268_r;
    reg node268_l;
    reg node269_r;
    reg node269_l;
    reg node270;
    reg node271;
    reg node272_r;
    reg node272_l;
    reg node273;
    reg node274;
    reg node275;
    reg node276_r;
    reg node276_l;
    reg node277_r;
    reg node277_l;
    reg node278_r;
    reg node278_l;
    reg node279_r;
    reg node279_l;
    reg node280;
    reg node281;
    reg node282;
    reg node283_r;
    reg node283_l;
    reg node284_r;
    reg node284_l;
    reg node285;
    reg node286;
    reg node287_r;
    reg node287_l;
    reg node288;
    reg node289;
    reg node290;
    reg node291_r;
    reg node291_l;
    reg node292_r;
    reg node292_l;
    reg node293_r;
    reg node293_l;
    reg node294_r;
    reg node294_l;
    reg node295_r;
    reg node295_l;
    reg node296;
    reg node297;
    reg node298_r;
    reg node298_l;
    reg node299;
    reg node300;
    reg node301_r;
    reg node301_l;
    reg node302_r;
    reg node302_l;
    reg node303;
    reg node304;
    reg node305_r;
    reg node305_l;
    reg node306;
    reg node307;
    reg node308_r;
    reg node308_l;
    reg node309_r;
    reg node309_l;
    reg node310_r;
    reg node310_l;
    reg node311;
    reg node312;
    reg node313_r;
    reg node313_l;
    reg node314;
    reg node315;
    reg node316_r;
    reg node316_l;
    reg node317_r;
    reg node317_l;
    reg node318;
    reg node319;
    reg node320_r;
    reg node320_l;
    reg node321;
    reg node322;
    reg node323_r;
    reg node323_l;
    reg node324_r;
    reg node324_l;
    reg node325_r;
    reg node325_l;
    reg node326_r;
    reg node326_l;
    reg node327;
    reg node328;
    reg node329_r;
    reg node329_l;
    reg node330;
    reg node331;
    reg node332_r;
    reg node332_l;
    reg node333_r;
    reg node333_l;
    reg node334;
    reg node335;
    reg node336_r;
    reg node336_l;
    reg node337;
    reg node338;
    reg node339_r;
    reg node339_l;
    reg node340_r;
    reg node340_l;
    reg node341_r;
    reg node341_l;
    reg node342;
    reg node343;
    reg node344_r;
    reg node344_l;
    reg node345;
    reg node346;
    reg node347_r;
    reg node347_l;
    reg node348_r;
    reg node348_l;
    reg node349;
    reg node350;
    reg node351_r;
    reg node351_l;
    reg node352;
    reg node353;
    reg node354_r;
    reg node354_l;
    reg node355_r;
    reg node355_l;
    reg node356_r;
    reg node356_l;
    reg node357_r;
    reg node357_l;
    reg node358_r;
    reg node358_l;
    reg node359_r;
    reg node359_l;
    reg node360;
    reg node361;
    reg node362_r;
    reg node362_l;
    reg node363;
    reg node364;
    reg node365_r;
    reg node365_l;
    reg node366_r;
    reg node366_l;
    reg node367;
    reg node368;
    reg node369_r;
    reg node369_l;
    reg node370;
    reg node371;
    reg node372_r;
    reg node372_l;
    reg node373_r;
    reg node373_l;
    reg node374_r;
    reg node374_l;
    reg node375;
    reg node376;
    reg node377_r;
    reg node377_l;
    reg node378;
    reg node379;
    reg node380_r;
    reg node380_l;
    reg node381_r;
    reg node381_l;
    reg node382;
    reg node383;
    reg node384_r;
    reg node384_l;
    reg node385;
    reg node386;
    reg node387_r;
    reg node387_l;
    reg node388_r;
    reg node388_l;
    reg node389_r;
    reg node389_l;
    reg node390_r;
    reg node390_l;
    reg node391;
    reg node392;
    reg node393;
    reg node394_r;
    reg node394_l;
    reg node395_r;
    reg node395_l;
    reg node396;
    reg node397;
    reg node398;
    reg node399_r;
    reg node399_l;
    reg node400_r;
    reg node400_l;
    reg node401;
    reg node402;
    reg node403_r;
    reg node403_l;
    reg node404_r;
    reg node404_l;
    reg node405;
    reg node406;
    reg node407_r;
    reg node407_l;
    reg node408;
    reg node409;
    reg node410;
    reg node411_r;
    reg node411_l;
    reg node412_r;
    reg node412_l;
    reg node413_r;
    reg node413_l;
    reg node414_r;
    reg node414_l;
    reg node415_r;
    reg node415_l;
    reg node416_r;
    reg node416_l;
    reg node417_r;
    reg node417_l;
    reg node418_r;
    reg node418_l;
    reg node419;
    reg node420;
    reg node421_r;
    reg node421_l;
    reg node422;
    reg node423;
    reg node424_r;
    reg node424_l;
    reg node425_r;
    reg node425_l;
    reg node426;
    reg node427;
    reg node428_r;
    reg node428_l;
    reg node429;
    reg node430;
    reg node431_r;
    reg node431_l;
    reg node432_r;
    reg node432_l;
    reg node433_r;
    reg node433_l;
    reg node434;
    reg node435;
    reg node436_r;
    reg node436_l;
    reg node437;
    reg node438;
    reg node439;
    reg node440_r;
    reg node440_l;
    reg node441_r;
    reg node441_l;
    reg node442_r;
    reg node442_l;
    reg node443_r;
    reg node443_l;
    reg node444;
    reg node445;
    reg node446_r;
    reg node446_l;
    reg node447;
    reg node448;
    reg node449_r;
    reg node449_l;
    reg node450_r;
    reg node450_l;
    reg node451;
    reg node452;
    reg node453_r;
    reg node453_l;
    reg node454;
    reg node455;
    reg node456_r;
    reg node456_l;
    reg node457_r;
    reg node457_l;
    reg node458_r;
    reg node458_l;
    reg node459;
    reg node460;
    reg node461;
    reg node462_r;
    reg node462_l;
    reg node463_r;
    reg node463_l;
    reg node464;
    reg node465;
    reg node466_r;
    reg node466_l;
    reg node467;
    reg node468;
    reg node469_r;
    reg node469_l;
    reg node470_r;
    reg node470_l;
    reg node471_r;
    reg node471_l;
    reg node472_r;
    reg node472_l;
    reg node473_r;
    reg node473_l;
    reg node474;
    reg node475;
    reg node476_r;
    reg node476_l;
    reg node477;
    reg node478;
    reg node479_r;
    reg node479_l;
    reg node480_r;
    reg node480_l;
    reg node481;
    reg node482;
    reg node483;
    reg node484_r;
    reg node484_l;
    reg node485_r;
    reg node485_l;
    reg node486_r;
    reg node486_l;
    reg node487;
    reg node488;
    reg node489_r;
    reg node489_l;
    reg node490;
    reg node491;
    reg node492_r;
    reg node492_l;
    reg node493;
    reg node494_r;
    reg node494_l;
    reg node495;
    reg node496;
    reg node497_r;
    reg node497_l;
    reg node498_r;
    reg node498_l;
    reg node499_r;
    reg node499_l;
    reg node500_r;
    reg node500_l;
    reg node501;
    reg node502;
    reg node503_r;
    reg node503_l;
    reg node504;
    reg node505;
    reg node506;
    reg node507_r;
    reg node507_l;
    reg node508_r;
    reg node508_l;
    reg node509;
    reg node510;
    reg node511_r;
    reg node511_l;
    reg node512_r;
    reg node512_l;
    reg node513;
    reg node514;
    reg node515_r;
    reg node515_l;
    reg node516;
    reg node517;
    reg node518_r;
    reg node518_l;
    reg node519_r;
    reg node519_l;
    reg node520_r;
    reg node520_l;
    reg node521_r;
    reg node521_l;
    reg node522_r;
    reg node522_l;
    reg node523_r;
    reg node523_l;
    reg node524;
    reg node525;
    reg node526_r;
    reg node526_l;
    reg node527;
    reg node528;
    reg node529_r;
    reg node529_l;
    reg node530_r;
    reg node530_l;
    reg node531;
    reg node532;
    reg node533;
    reg node534_r;
    reg node534_l;
    reg node535_r;
    reg node535_l;
    reg node536_r;
    reg node536_l;
    reg node537;
    reg node538;
    reg node539_r;
    reg node539_l;
    reg node540;
    reg node541;
    reg node542_r;
    reg node542_l;
    reg node543_r;
    reg node543_l;
    reg node544;
    reg node545;
    reg node546_r;
    reg node546_l;
    reg node547;
    reg node548;
    reg node549_r;
    reg node549_l;
    reg node550_r;
    reg node550_l;
    reg node551_r;
    reg node551_l;
    reg node552_r;
    reg node552_l;
    reg node553;
    reg node554;
    reg node555_r;
    reg node555_l;
    reg node556;
    reg node557;
    reg node558_r;
    reg node558_l;
    reg node559_r;
    reg node559_l;
    reg node560;
    reg node561;
    reg node562_r;
    reg node562_l;
    reg node563;
    reg node564;
    reg node565_r;
    reg node565_l;
    reg node566_r;
    reg node566_l;
    reg node567_r;
    reg node567_l;
    reg node568;
    reg node569;
    reg node570_r;
    reg node570_l;
    reg node571;
    reg node572;
    reg node573_r;
    reg node573_l;
    reg node574_r;
    reg node574_l;
    reg node575;
    reg node576;
    reg node577_r;
    reg node577_l;
    reg node578;
    reg node579;
    reg node580_r;
    reg node580_l;
    reg node581_r;
    reg node581_l;
    reg node582_r;
    reg node582_l;
    reg node583_r;
    reg node583_l;
    reg node584_r;
    reg node584_l;
    reg node585;
    reg node586;
    reg node587_r;
    reg node587_l;
    reg node588;
    reg node589;
    reg node590_r;
    reg node590_l;
    reg node591_r;
    reg node591_l;
    reg node592;
    reg node593;
    reg node594_r;
    reg node594_l;
    reg node595;
    reg node596;
    reg node597_r;
    reg node597_l;
    reg node598_r;
    reg node598_l;
    reg node599_r;
    reg node599_l;
    reg node600;
    reg node601;
    reg node602_r;
    reg node602_l;
    reg node603;
    reg node604;
    reg node605_r;
    reg node605_l;
    reg node606_r;
    reg node606_l;
    reg node607;
    reg node608;
    reg node609_r;
    reg node609_l;
    reg node610;
    reg node611;
    reg node612_r;
    reg node612_l;
    reg node613_r;
    reg node613_l;
    reg node614_r;
    reg node614_l;
    reg node615_r;
    reg node615_l;
    reg node616;
    reg node617;
    reg node618_r;
    reg node618_l;
    reg node619;
    reg node620;
    reg node621_r;
    reg node621_l;
    reg node622_r;
    reg node622_l;
    reg node623;
    reg node624;
    reg node625_r;
    reg node625_l;
    reg node626;
    reg node627;
    reg node628_r;
    reg node628_l;
    reg node629_r;
    reg node629_l;
    reg node630_r;
    reg node630_l;
    reg node631;
    reg node632;
    reg node633_r;
    reg node633_l;
    reg node634;
    reg node635;
    reg node636_r;
    reg node636_l;
    reg node637_r;
    reg node637_l;
    reg node638;
    reg node639;
    reg node640_r;
    reg node640_l;
    reg node641;
    reg node642;
    reg node643_r;
    reg node643_l;
    reg node644_r;
    reg node644_l;
    reg node645_r;
    reg node645_l;
    reg node646_r;
    reg node646_l;
    reg node647_r;
    reg node647_l;
    reg node648_r;
    reg node648_l;
    reg node649_r;
    reg node649_l;
    reg node650;
    reg node651;
    reg node652_r;
    reg node652_l;
    reg node653;
    reg node654;
    reg node655_r;
    reg node655_l;
    reg node656_r;
    reg node656_l;
    reg node657;
    reg node658;
    reg node659_r;
    reg node659_l;
    reg node660;
    reg node661;
    reg node662_r;
    reg node662_l;
    reg node663_r;
    reg node663_l;
    reg node664;
    reg node665_r;
    reg node665_l;
    reg node666;
    reg node667;
    reg node668_r;
    reg node668_l;
    reg node669_r;
    reg node669_l;
    reg node670;
    reg node671;
    reg node672;
    reg node673_r;
    reg node673_l;
    reg node674_r;
    reg node674_l;
    reg node675_r;
    reg node675_l;
    reg node676_r;
    reg node676_l;
    reg node677;
    reg node678;
    reg node679_r;
    reg node679_l;
    reg node680;
    reg node681;
    reg node682_r;
    reg node682_l;
    reg node683_r;
    reg node683_l;
    reg node684;
    reg node685;
    reg node686_r;
    reg node686_l;
    reg node687;
    reg node688;
    reg node689_r;
    reg node689_l;
    reg node690_r;
    reg node690_l;
    reg node691_r;
    reg node691_l;
    reg node692;
    reg node693;
    reg node694_r;
    reg node694_l;
    reg node695;
    reg node696;
    reg node697_r;
    reg node697_l;
    reg node698_r;
    reg node698_l;
    reg node699;
    reg node700;
    reg node701_r;
    reg node701_l;
    reg node702;
    reg node703;
    reg node704_r;
    reg node704_l;
    reg node705_r;
    reg node705_l;
    reg node706_r;
    reg node706_l;
    reg node707_r;
    reg node707_l;
    reg node708_r;
    reg node708_l;
    reg node709;
    reg node710;
    reg node711_r;
    reg node711_l;
    reg node712;
    reg node713;
    reg node714_r;
    reg node714_l;
    reg node715_r;
    reg node715_l;
    reg node716;
    reg node717;
    reg node718_r;
    reg node718_l;
    reg node719;
    reg node720;
    reg node721_r;
    reg node721_l;
    reg node722_r;
    reg node722_l;
    reg node723_r;
    reg node723_l;
    reg node724;
    reg node725;
    reg node726_r;
    reg node726_l;
    reg node727;
    reg node728;
    reg node729_r;
    reg node729_l;
    reg node730_r;
    reg node730_l;
    reg node731;
    reg node732;
    reg node733_r;
    reg node733_l;
    reg node734;
    reg node735;
    reg node736_r;
    reg node736_l;
    reg node737_r;
    reg node737_l;
    reg node738_r;
    reg node738_l;
    reg node739_r;
    reg node739_l;
    reg node740;
    reg node741;
    reg node742_r;
    reg node742_l;
    reg node743;
    reg node744;
    reg node745_r;
    reg node745_l;
    reg node746_r;
    reg node746_l;
    reg node747;
    reg node748;
    reg node749_r;
    reg node749_l;
    reg node750;
    reg node751;
    reg node752_r;
    reg node752_l;
    reg node753_r;
    reg node753_l;
    reg node754_r;
    reg node754_l;
    reg node755;
    reg node756;
    reg node757_r;
    reg node757_l;
    reg node758;
    reg node759;
    reg node760_r;
    reg node760_l;
    reg node761_r;
    reg node761_l;
    reg node762;
    reg node763;
    reg node764_r;
    reg node764_l;
    reg node765;
    reg node766;
    reg node767_r;
    reg node767_l;
    reg node768_r;
    reg node768_l;
    reg node769_r;
    reg node769_l;
    reg node770_r;
    reg node770_l;
    reg node771_r;
    reg node771_l;
    reg node772_r;
    reg node772_l;
    reg node773;
    reg node774;
    reg node775_r;
    reg node775_l;
    reg node776;
    reg node777;
    reg node778_r;
    reg node778_l;
    reg node779_r;
    reg node779_l;
    reg node780;
    reg node781;
    reg node782_r;
    reg node782_l;
    reg node783;
    reg node784;
    reg node785;
    reg node786_r;
    reg node786_l;
    reg node787_r;
    reg node787_l;
    reg node788_r;
    reg node788_l;
    reg node789_r;
    reg node789_l;
    reg node790;
    reg node791;
    reg node792_r;
    reg node792_l;
    reg node793;
    reg node794;
    reg node795_r;
    reg node795_l;
    reg node796_r;
    reg node796_l;
    reg node797;
    reg node798;
    reg node799_r;
    reg node799_l;
    reg node800;
    reg node801;
    reg node802_r;
    reg node802_l;
    reg node803_r;
    reg node803_l;
    reg node804_r;
    reg node804_l;
    reg node805;
    reg node806;
    reg node807_r;
    reg node807_l;
    reg node808;
    reg node809;
    reg node810_r;
    reg node810_l;
    reg node811_r;
    reg node811_l;
    reg node812;
    reg node813;
    reg node814;
    reg node815_r;
    reg node815_l;
    reg node816_r;
    reg node816_l;
    reg node817_r;
    reg node817_l;
    reg node818_r;
    reg node818_l;
    reg node819_r;
    reg node819_l;
    reg node820;
    reg node821;
    reg node822;
    reg node823_r;
    reg node823_l;
    reg node824_r;
    reg node824_l;
    reg node825;
    reg node826;
    reg node827_r;
    reg node827_l;
    reg node828;
    reg node829;
    reg node830_r;
    reg node830_l;
    reg node831_r;
    reg node831_l;
    reg node832;
    reg node833;
    reg node834;
    reg node835_r;
    reg node835_l;
    reg node836_r;
    reg node836_l;
    reg node837_r;
    reg node837_l;
    reg node838;
    reg node839_r;
    reg node839_l;
    reg node840;
    reg node841;
    reg node842_r;
    reg node842_l;
    reg node843;
    reg node844_r;
    reg node844_l;
    reg node845;
    reg node846;
    reg node847_r;
    reg node847_l;
    reg node848_r;
    reg node848_l;
    reg node849;
    reg node850_r;
    reg node850_l;
    reg node851;
    reg node852;
    reg node853_r;
    reg node853_l;
    reg node854;
    reg node855_r;
    reg node855_l;
    reg node856;
    reg node857;
    reg node858_r;
    reg node858_l;
    reg node859_r;
    reg node859_l;
    reg node860_r;
    reg node860_l;
    reg node861_r;
    reg node861_l;
    reg node862_r;
    reg node862_l;
    reg node863_r;
    reg node863_l;
    reg node864_r;
    reg node864_l;
    reg node865_r;
    reg node865_l;
    reg node866_r;
    reg node866_l;
    reg node867;
    reg node868;
    reg node869_r;
    reg node869_l;
    reg node870;
    reg node871;
    reg node872_r;
    reg node872_l;
    reg node873_r;
    reg node873_l;
    reg node874;
    reg node875;
    reg node876_r;
    reg node876_l;
    reg node877;
    reg node878;
    reg node879_r;
    reg node879_l;
    reg node880_r;
    reg node880_l;
    reg node881_r;
    reg node881_l;
    reg node882;
    reg node883;
    reg node884_r;
    reg node884_l;
    reg node885;
    reg node886;
    reg node887_r;
    reg node887_l;
    reg node888_r;
    reg node888_l;
    reg node889;
    reg node890;
    reg node891_r;
    reg node891_l;
    reg node892;
    reg node893;
    reg node894_r;
    reg node894_l;
    reg node895_r;
    reg node895_l;
    reg node896_r;
    reg node896_l;
    reg node897_r;
    reg node897_l;
    reg node898;
    reg node899;
    reg node900_r;
    reg node900_l;
    reg node901;
    reg node902;
    reg node903_r;
    reg node903_l;
    reg node904_r;
    reg node904_l;
    reg node905;
    reg node906;
    reg node907;
    reg node908_r;
    reg node908_l;
    reg node909_r;
    reg node909_l;
    reg node910_r;
    reg node910_l;
    reg node911;
    reg node912;
    reg node913_r;
    reg node913_l;
    reg node914;
    reg node915;
    reg node916_r;
    reg node916_l;
    reg node917_r;
    reg node917_l;
    reg node918;
    reg node919;
    reg node920_r;
    reg node920_l;
    reg node921;
    reg node922;
    reg node923_r;
    reg node923_l;
    reg node924_r;
    reg node924_l;
    reg node925_r;
    reg node925_l;
    reg node926_r;
    reg node926_l;
    reg node927_r;
    reg node927_l;
    reg node928;
    reg node929;
    reg node930_r;
    reg node930_l;
    reg node931;
    reg node932;
    reg node933_r;
    reg node933_l;
    reg node934_r;
    reg node934_l;
    reg node935;
    reg node936;
    reg node937_r;
    reg node937_l;
    reg node938;
    reg node939;
    reg node940_r;
    reg node940_l;
    reg node941;
    reg node942;
    reg node943_r;
    reg node943_l;
    reg node944_r;
    reg node944_l;
    reg node945_r;
    reg node945_l;
    reg node946_r;
    reg node946_l;
    reg node947;
    reg node948;
    reg node949_r;
    reg node949_l;
    reg node950;
    reg node951;
    reg node952_r;
    reg node952_l;
    reg node953_r;
    reg node953_l;
    reg node954;
    reg node955;
    reg node956_r;
    reg node956_l;
    reg node957;
    reg node958;
    reg node959_r;
    reg node959_l;
    reg node960_r;
    reg node960_l;
    reg node961_r;
    reg node961_l;
    reg node962;
    reg node963;
    reg node964_r;
    reg node964_l;
    reg node965;
    reg node966;
    reg node967_r;
    reg node967_l;
    reg node968_r;
    reg node968_l;
    reg node969;
    reg node970;
    reg node971_r;
    reg node971_l;
    reg node972;
    reg node973;
    reg node974_r;
    reg node974_l;
    reg node975_r;
    reg node975_l;
    reg node976_r;
    reg node976_l;
    reg node977_r;
    reg node977_l;
    reg node978_r;
    reg node978_l;
    reg node979_r;
    reg node979_l;
    reg node980;
    reg node981;
    reg node982_r;
    reg node982_l;
    reg node983;
    reg node984;
    reg node985_r;
    reg node985_l;
    reg node986_r;
    reg node986_l;
    reg node987;
    reg node988;
    reg node989;
    reg node990_r;
    reg node990_l;
    reg node991_r;
    reg node991_l;
    reg node992_r;
    reg node992_l;
    reg node993;
    reg node994;
    reg node995;
    reg node996_r;
    reg node996_l;
    reg node997_r;
    reg node997_l;
    reg node998;
    reg node999;
    reg node1000;
    reg node1001_r;
    reg node1001_l;
    reg node1002_r;
    reg node1002_l;
    reg node1003_r;
    reg node1003_l;
    reg node1004_r;
    reg node1004_l;
    reg node1005;
    reg node1006;
    reg node1007_r;
    reg node1007_l;
    reg node1008;
    reg node1009;
    reg node1010_r;
    reg node1010_l;
    reg node1011_r;
    reg node1011_l;
    reg node1012;
    reg node1013;
    reg node1014_r;
    reg node1014_l;
    reg node1015;
    reg node1016;
    reg node1017_r;
    reg node1017_l;
    reg node1018_r;
    reg node1018_l;
    reg node1019_r;
    reg node1019_l;
    reg node1020;
    reg node1021;
    reg node1022_r;
    reg node1022_l;
    reg node1023;
    reg node1024;
    reg node1025_r;
    reg node1025_l;
    reg node1026_r;
    reg node1026_l;
    reg node1027;
    reg node1028;
    reg node1029_r;
    reg node1029_l;
    reg node1030;
    reg node1031;
    reg node1032_r;
    reg node1032_l;
    reg node1033_r;
    reg node1033_l;
    reg node1034_r;
    reg node1034_l;
    reg node1035_r;
    reg node1035_l;
    reg node1036_r;
    reg node1036_l;
    reg node1037;
    reg node1038;
    reg node1039_r;
    reg node1039_l;
    reg node1040;
    reg node1041;
    reg node1042_r;
    reg node1042_l;
    reg node1043_r;
    reg node1043_l;
    reg node1044;
    reg node1045;
    reg node1046_r;
    reg node1046_l;
    reg node1047;
    reg node1048;
    reg node1049_r;
    reg node1049_l;
    reg node1050_r;
    reg node1050_l;
    reg node1051_r;
    reg node1051_l;
    reg node1052;
    reg node1053;
    reg node1054_r;
    reg node1054_l;
    reg node1055;
    reg node1056;
    reg node1057_r;
    reg node1057_l;
    reg node1058_r;
    reg node1058_l;
    reg node1059;
    reg node1060;
    reg node1061_r;
    reg node1061_l;
    reg node1062;
    reg node1063;
    reg node1064_r;
    reg node1064_l;
    reg node1065_r;
    reg node1065_l;
    reg node1066_r;
    reg node1066_l;
    reg node1067_r;
    reg node1067_l;
    reg node1068;
    reg node1069;
    reg node1070_r;
    reg node1070_l;
    reg node1071;
    reg node1072;
    reg node1073_r;
    reg node1073_l;
    reg node1074_r;
    reg node1074_l;
    reg node1075;
    reg node1076;
    reg node1077_r;
    reg node1077_l;
    reg node1078;
    reg node1079;
    reg node1080_r;
    reg node1080_l;
    reg node1081_r;
    reg node1081_l;
    reg node1082_r;
    reg node1082_l;
    reg node1083;
    reg node1084;
    reg node1085_r;
    reg node1085_l;
    reg node1086;
    reg node1087;
    reg node1088_r;
    reg node1088_l;
    reg node1089_r;
    reg node1089_l;
    reg node1090;
    reg node1091;
    reg node1092_r;
    reg node1092_l;
    reg node1093;
    reg node1094;
    reg node1095_r;
    reg node1095_l;
    reg node1096_r;
    reg node1096_l;
    reg node1097_r;
    reg node1097_l;
    reg node1098_r;
    reg node1098_l;
    reg node1099_r;
    reg node1099_l;
    reg node1100_r;
    reg node1100_l;
    reg node1101_r;
    reg node1101_l;
    reg node1102;
    reg node1103;
    reg node1104_r;
    reg node1104_l;
    reg node1105;
    reg node1106;
    reg node1107_r;
    reg node1107_l;
    reg node1108_r;
    reg node1108_l;
    reg node1109;
    reg node1110;
    reg node1111_r;
    reg node1111_l;
    reg node1112;
    reg node1113;
    reg node1114_r;
    reg node1114_l;
    reg node1115_r;
    reg node1115_l;
    reg node1116_r;
    reg node1116_l;
    reg node1117;
    reg node1118;
    reg node1119_r;
    reg node1119_l;
    reg node1120;
    reg node1121;
    reg node1122_r;
    reg node1122_l;
    reg node1123_r;
    reg node1123_l;
    reg node1124;
    reg node1125;
    reg node1126_r;
    reg node1126_l;
    reg node1127;
    reg node1128;
    reg node1129_r;
    reg node1129_l;
    reg node1130_r;
    reg node1130_l;
    reg node1131_r;
    reg node1131_l;
    reg node1132_r;
    reg node1132_l;
    reg node1133;
    reg node1134;
    reg node1135_r;
    reg node1135_l;
    reg node1136;
    reg node1137;
    reg node1138_r;
    reg node1138_l;
    reg node1139_r;
    reg node1139_l;
    reg node1140;
    reg node1141;
    reg node1142_r;
    reg node1142_l;
    reg node1143;
    reg node1144;
    reg node1145_r;
    reg node1145_l;
    reg node1146_r;
    reg node1146_l;
    reg node1147_r;
    reg node1147_l;
    reg node1148;
    reg node1149;
    reg node1150_r;
    reg node1150_l;
    reg node1151;
    reg node1152;
    reg node1153_r;
    reg node1153_l;
    reg node1154_r;
    reg node1154_l;
    reg node1155;
    reg node1156;
    reg node1157_r;
    reg node1157_l;
    reg node1158;
    reg node1159;
    reg node1160_r;
    reg node1160_l;
    reg node1161_r;
    reg node1161_l;
    reg node1162_r;
    reg node1162_l;
    reg node1163_r;
    reg node1163_l;
    reg node1164_r;
    reg node1164_l;
    reg node1165;
    reg node1166;
    reg node1167;
    reg node1168;
    reg node1169_r;
    reg node1169_l;
    reg node1170_r;
    reg node1170_l;
    reg node1171_r;
    reg node1171_l;
    reg node1172;
    reg node1173;
    reg node1174_r;
    reg node1174_l;
    reg node1175;
    reg node1176;
    reg node1177_r;
    reg node1177_l;
    reg node1178_r;
    reg node1178_l;
    reg node1179;
    reg node1180;
    reg node1181;
    reg node1182_r;
    reg node1182_l;
    reg node1183_r;
    reg node1183_l;
    reg node1184_r;
    reg node1184_l;
    reg node1185_r;
    reg node1185_l;
    reg node1186;
    reg node1187;
    reg node1188_r;
    reg node1188_l;
    reg node1189;
    reg node1190;
    reg node1191_r;
    reg node1191_l;
    reg node1192_r;
    reg node1192_l;
    reg node1193;
    reg node1194;
    reg node1195_r;
    reg node1195_l;
    reg node1196;
    reg node1197;
    reg node1198_r;
    reg node1198_l;
    reg node1199_r;
    reg node1199_l;
    reg node1200_r;
    reg node1200_l;
    reg node1201;
    reg node1202;
    reg node1203;
    reg node1204_r;
    reg node1204_l;
    reg node1205_r;
    reg node1205_l;
    reg node1206;
    reg node1207;
    reg node1208_r;
    reg node1208_l;
    reg node1209;
    reg node1210;
    reg node1211_r;
    reg node1211_l;
    reg node1212_r;
    reg node1212_l;
    reg node1213_r;
    reg node1213_l;
    reg node1214_r;
    reg node1214_l;
    reg node1215_r;
    reg node1215_l;
    reg node1216_r;
    reg node1216_l;
    reg node1217;
    reg node1218;
    reg node1219_r;
    reg node1219_l;
    reg node1220;
    reg node1221;
    reg node1222_r;
    reg node1222_l;
    reg node1223_r;
    reg node1223_l;
    reg node1224;
    reg node1225;
    reg node1226_r;
    reg node1226_l;
    reg node1227;
    reg node1228;
    reg node1229;
    reg node1230;
    reg node1231_r;
    reg node1231_l;
    reg node1232_r;
    reg node1232_l;
    reg node1233_r;
    reg node1233_l;
    reg node1234_r;
    reg node1234_l;
    reg node1235;
    reg node1236;
    reg node1237;
    reg node1238_r;
    reg node1238_l;
    reg node1239_r;
    reg node1239_l;
    reg node1240_r;
    reg node1240_l;
    reg node1241;
    reg node1242;
    reg node1243_r;
    reg node1243_l;
    reg node1244;
    reg node1245;
    reg node1246_r;
    reg node1246_l;
    reg node1247_r;
    reg node1247_l;
    reg node1248;
    reg node1249;
    reg node1250;
    reg node1251_r;
    reg node1251_l;
    reg node1252_r;
    reg node1252_l;
    reg node1253;
    reg node1254;
    reg node1255_r;
    reg node1255_l;
    reg node1256_r;
    reg node1256_l;
    reg node1257;
    reg node1258;
    reg node1259_r;
    reg node1259_l;
    reg node1260;
    reg node1261;
    reg node1262_r;
    reg node1262_l;
    reg node1263_r;
    reg node1263_l;
    reg node1264_r;
    reg node1264_l;
    reg node1265_r;
    reg node1265_l;
    reg node1266_r;
    reg node1266_l;
    reg node1267_r;
    reg node1267_l;
    reg node1268_r;
    reg node1268_l;
    reg node1269_r;
    reg node1269_l;
    reg node1270;
    reg node1271;
    reg node1272_r;
    reg node1272_l;
    reg node1273;
    reg node1274;
    reg node1275_r;
    reg node1275_l;
    reg node1276_r;
    reg node1276_l;
    reg node1277;
    reg node1278;
    reg node1279_r;
    reg node1279_l;
    reg node1280;
    reg node1281;
    reg node1282_r;
    reg node1282_l;
    reg node1283_r;
    reg node1283_l;
    reg node1284_r;
    reg node1284_l;
    reg node1285;
    reg node1286;
    reg node1287_r;
    reg node1287_l;
    reg node1288;
    reg node1289;
    reg node1290_r;
    reg node1290_l;
    reg node1291_r;
    reg node1291_l;
    reg node1292;
    reg node1293;
    reg node1294_r;
    reg node1294_l;
    reg node1295;
    reg node1296;
    reg node1297_r;
    reg node1297_l;
    reg node1298_r;
    reg node1298_l;
    reg node1299_r;
    reg node1299_l;
    reg node1300_r;
    reg node1300_l;
    reg node1301;
    reg node1302;
    reg node1303_r;
    reg node1303_l;
    reg node1304;
    reg node1305;
    reg node1306_r;
    reg node1306_l;
    reg node1307_r;
    reg node1307_l;
    reg node1308;
    reg node1309;
    reg node1310_r;
    reg node1310_l;
    reg node1311;
    reg node1312;
    reg node1313_r;
    reg node1313_l;
    reg node1314_r;
    reg node1314_l;
    reg node1315_r;
    reg node1315_l;
    reg node1316;
    reg node1317;
    reg node1318_r;
    reg node1318_l;
    reg node1319;
    reg node1320;
    reg node1321_r;
    reg node1321_l;
    reg node1322_r;
    reg node1322_l;
    reg node1323;
    reg node1324;
    reg node1325;
    reg node1326_r;
    reg node1326_l;
    reg node1327_r;
    reg node1327_l;
    reg node1328_r;
    reg node1328_l;
    reg node1329_r;
    reg node1329_l;
    reg node1330_r;
    reg node1330_l;
    reg node1331;
    reg node1332;
    reg node1333_r;
    reg node1333_l;
    reg node1334;
    reg node1335;
    reg node1336;
    reg node1337_r;
    reg node1337_l;
    reg node1338_r;
    reg node1338_l;
    reg node1339_r;
    reg node1339_l;
    reg node1340;
    reg node1341;
    reg node1342_r;
    reg node1342_l;
    reg node1343;
    reg node1344;
    reg node1345_r;
    reg node1345_l;
    reg node1346_r;
    reg node1346_l;
    reg node1347;
    reg node1348;
    reg node1349_r;
    reg node1349_l;
    reg node1350;
    reg node1351;
    reg node1352_r;
    reg node1352_l;
    reg node1353_r;
    reg node1353_l;
    reg node1354_r;
    reg node1354_l;
    reg node1355_r;
    reg node1355_l;
    reg node1356;
    reg node1357;
    reg node1358_r;
    reg node1358_l;
    reg node1359;
    reg node1360;
    reg node1361_r;
    reg node1361_l;
    reg node1362_r;
    reg node1362_l;
    reg node1363;
    reg node1364;
    reg node1365_r;
    reg node1365_l;
    reg node1366;
    reg node1367;
    reg node1368_r;
    reg node1368_l;
    reg node1369_r;
    reg node1369_l;
    reg node1370;
    reg node1371;
    reg node1372_r;
    reg node1372_l;
    reg node1373_r;
    reg node1373_l;
    reg node1374;
    reg node1375;
    reg node1376_r;
    reg node1376_l;
    reg node1377;
    reg node1378;
    reg node1379_r;
    reg node1379_l;
    reg node1380_r;
    reg node1380_l;
    reg node1381_r;
    reg node1381_l;
    reg node1382_r;
    reg node1382_l;
    reg node1383_r;
    reg node1383_l;
    reg node1384_r;
    reg node1384_l;
    reg node1385;
    reg node1386;
    reg node1387_r;
    reg node1387_l;
    reg node1388;
    reg node1389;
    reg node1390_r;
    reg node1390_l;
    reg node1391_r;
    reg node1391_l;
    reg node1392;
    reg node1393;
    reg node1394_r;
    reg node1394_l;
    reg node1395;
    reg node1396;
    reg node1397_r;
    reg node1397_l;
    reg node1398_r;
    reg node1398_l;
    reg node1399_r;
    reg node1399_l;
    reg node1400;
    reg node1401;
    reg node1402;
    reg node1403_r;
    reg node1403_l;
    reg node1404_r;
    reg node1404_l;
    reg node1405;
    reg node1406;
    reg node1407_r;
    reg node1407_l;
    reg node1408;
    reg node1409;
    reg node1410_r;
    reg node1410_l;
    reg node1411_r;
    reg node1411_l;
    reg node1412_r;
    reg node1412_l;
    reg node1413_r;
    reg node1413_l;
    reg node1414;
    reg node1415;
    reg node1416_r;
    reg node1416_l;
    reg node1417;
    reg node1418;
    reg node1419;
    reg node1420_r;
    reg node1420_l;
    reg node1421;
    reg node1422;
    reg node1423_r;
    reg node1423_l;
    reg node1424_r;
    reg node1424_l;
    reg node1425_r;
    reg node1425_l;
    reg node1426_r;
    reg node1426_l;
    reg node1427_r;
    reg node1427_l;
    reg node1428;
    reg node1429;
    reg node1430_r;
    reg node1430_l;
    reg node1431;
    reg node1432;
    reg node1433_r;
    reg node1433_l;
    reg node1434_r;
    reg node1434_l;
    reg node1435;
    reg node1436;
    reg node1437_r;
    reg node1437_l;
    reg node1438;
    reg node1439;
    reg node1440_r;
    reg node1440_l;
    reg node1441_r;
    reg node1441_l;
    reg node1442_r;
    reg node1442_l;
    reg node1443;
    reg node1444;
    reg node1445;
    reg node1446_r;
    reg node1446_l;
    reg node1447_r;
    reg node1447_l;
    reg node1448;
    reg node1449;
    reg node1450_r;
    reg node1450_l;
    reg node1451;
    reg node1452;
    reg node1453_r;
    reg node1453_l;
    reg node1454_r;
    reg node1454_l;
    reg node1455_r;
    reg node1455_l;
    reg node1456;
    reg node1457;
    reg node1458_r;
    reg node1458_l;
    reg node1459;
    reg node1460_r;
    reg node1460_l;
    reg node1461;
    reg node1462;
    reg node1463;
    reg node1464_r;
    reg node1464_l;
    reg node1465_r;
    reg node1465_l;
    reg node1466_r;
    reg node1466_l;
    reg node1467_r;
    reg node1467_l;
    reg node1468_r;
    reg node1468_l;
    reg node1469_r;
    reg node1469_l;
    reg node1470_r;
    reg node1470_l;
    reg node1471;
    reg node1472;
    reg node1473_r;
    reg node1473_l;
    reg node1474;
    reg node1475;
    reg node1476;
    reg node1477_r;
    reg node1477_l;
    reg node1478_r;
    reg node1478_l;
    reg node1479_r;
    reg node1479_l;
    reg node1480;
    reg node1481;
    reg node1482_r;
    reg node1482_l;
    reg node1483;
    reg node1484;
    reg node1485_r;
    reg node1485_l;
    reg node1486_r;
    reg node1486_l;
    reg node1487;
    reg node1488;
    reg node1489_r;
    reg node1489_l;
    reg node1490;
    reg node1491;
    reg node1492_r;
    reg node1492_l;
    reg node1493_r;
    reg node1493_l;
    reg node1494_r;
    reg node1494_l;
    reg node1495_r;
    reg node1495_l;
    reg node1496;
    reg node1497;
    reg node1498;
    reg node1499_r;
    reg node1499_l;
    reg node1500_r;
    reg node1500_l;
    reg node1501;
    reg node1502;
    reg node1503_r;
    reg node1503_l;
    reg node1504;
    reg node1505;
    reg node1506_r;
    reg node1506_l;
    reg node1507_r;
    reg node1507_l;
    reg node1508_r;
    reg node1508_l;
    reg node1509;
    reg node1510;
    reg node1511;
    reg node1512_r;
    reg node1512_l;
    reg node1513;
    reg node1514_r;
    reg node1514_l;
    reg node1515;
    reg node1516;
    reg node1517_r;
    reg node1517_l;
    reg node1518_r;
    reg node1518_l;
    reg node1519_r;
    reg node1519_l;
    reg node1520_r;
    reg node1520_l;
    reg node1521_r;
    reg node1521_l;
    reg node1522;
    reg node1523;
    reg node1524_r;
    reg node1524_l;
    reg node1525;
    reg node1526;
    reg node1527_r;
    reg node1527_l;
    reg node1528_r;
    reg node1528_l;
    reg node1529;
    reg node1530;
    reg node1531_r;
    reg node1531_l;
    reg node1532;
    reg node1533;
    reg node1534_r;
    reg node1534_l;
    reg node1535_r;
    reg node1535_l;
    reg node1536_r;
    reg node1536_l;
    reg node1537;
    reg node1538;
    reg node1539_r;
    reg node1539_l;
    reg node1540;
    reg node1541;
    reg node1542_r;
    reg node1542_l;
    reg node1543;
    reg node1544;
    reg node1545_r;
    reg node1545_l;
    reg node1546_r;
    reg node1546_l;
    reg node1547_r;
    reg node1547_l;
    reg node1548_r;
    reg node1548_l;
    reg node1549;
    reg node1550;
    reg node1551_r;
    reg node1551_l;
    reg node1552;
    reg node1553;
    reg node1554_r;
    reg node1554_l;
    reg node1555_r;
    reg node1555_l;
    reg node1556;
    reg node1557;
    reg node1558_r;
    reg node1558_l;
    reg node1559;
    reg node1560;
    reg node1561_r;
    reg node1561_l;
    reg node1562_r;
    reg node1562_l;
    reg node1563_r;
    reg node1563_l;
    reg node1564;
    reg node1565;
    reg node1566_r;
    reg node1566_l;
    reg node1567;
    reg node1568;
    reg node1569_r;
    reg node1569_l;
    reg node1570_r;
    reg node1570_l;
    reg node1571;
    reg node1572;
    reg node1573_r;
    reg node1573_l;
    reg node1574;
    reg node1575;
    reg node1576_r;
    reg node1576_l;
    reg node1577_r;
    reg node1577_l;
    reg node1578_r;
    reg node1578_l;
    reg node1579_r;
    reg node1579_l;
    reg node1580_r;
    reg node1580_l;
    reg node1581_r;
    reg node1581_l;
    reg node1582;
    reg node1583;
    reg node1584_r;
    reg node1584_l;
    reg node1585;
    reg node1586;
    reg node1587_r;
    reg node1587_l;
    reg node1588;
    reg node1589_r;
    reg node1589_l;
    reg node1590;
    reg node1591;
    reg node1592_r;
    reg node1592_l;
    reg node1593_r;
    reg node1593_l;
    reg node1594_r;
    reg node1594_l;
    reg node1595;
    reg node1596;
    reg node1597_r;
    reg node1597_l;
    reg node1598;
    reg node1599;
    reg node1600_r;
    reg node1600_l;
    reg node1601_r;
    reg node1601_l;
    reg node1602;
    reg node1603;
    reg node1604_r;
    reg node1604_l;
    reg node1605;
    reg node1606;
    reg node1607_r;
    reg node1607_l;
    reg node1608_r;
    reg node1608_l;
    reg node1609_r;
    reg node1609_l;
    reg node1610_r;
    reg node1610_l;
    reg node1611;
    reg node1612;
    reg node1613_r;
    reg node1613_l;
    reg node1614;
    reg node1615;
    reg node1616_r;
    reg node1616_l;
    reg node1617;
    reg node1618_r;
    reg node1618_l;
    reg node1619;
    reg node1620;
    reg node1621_r;
    reg node1621_l;
    reg node1622_r;
    reg node1622_l;
    reg node1623_r;
    reg node1623_l;
    reg node1624;
    reg node1625;
    reg node1626_r;
    reg node1626_l;
    reg node1627;
    reg node1628;
    reg node1629;
    reg node1630_r;
    reg node1630_l;
    reg node1631_r;
    reg node1631_l;
    reg node1632_r;
    reg node1632_l;
    reg node1633_r;
    reg node1633_l;
    reg node1634_r;
    reg node1634_l;
    reg node1635;
    reg node1636;
    reg node1637_r;
    reg node1637_l;
    reg node1638;
    reg node1639;
    reg node1640_r;
    reg node1640_l;
    reg node1641_r;
    reg node1641_l;
    reg node1642;
    reg node1643;
    reg node1644_r;
    reg node1644_l;
    reg node1645;
    reg node1646;
    reg node1647_r;
    reg node1647_l;
    reg node1648_r;
    reg node1648_l;
    reg node1649_r;
    reg node1649_l;
    reg node1650;
    reg node1651;
    reg node1652_r;
    reg node1652_l;
    reg node1653;
    reg node1654;
    reg node1655_r;
    reg node1655_l;
    reg node1656_r;
    reg node1656_l;
    reg node1657;
    reg node1658;
    reg node1659_r;
    reg node1659_l;
    reg node1660;
    reg node1661;
    reg node1662_r;
    reg node1662_l;
    reg node1663_r;
    reg node1663_l;
    reg node1664_r;
    reg node1664_l;
    reg node1665_r;
    reg node1665_l;
    reg node1666;
    reg node1667;
    reg node1668_r;
    reg node1668_l;
    reg node1669;
    reg node1670;
    reg node1671_r;
    reg node1671_l;
    reg node1672_r;
    reg node1672_l;
    reg node1673;
    reg node1674;
    reg node1675_r;
    reg node1675_l;
    reg node1676;
    reg node1677;
    reg node1678_r;
    reg node1678_l;
    reg node1679_r;
    reg node1679_l;
    reg node1680_r;
    reg node1680_l;
    reg node1681;
    reg node1682;
    reg node1683_r;
    reg node1683_l;
    reg node1684;
    reg node1685;
    reg node1686_r;
    reg node1686_l;
    reg node1687_r;
    reg node1687_l;
    reg node1688;
    reg node1689;
    reg node1690_r;
    reg node1690_l;
    reg node1691;
    reg node1692;
    reg result0;
    reg result1;
    reg result2;
    reg result3;
    reg result4;
    reg result5;
    reg result6;
    reg result7;
    reg result8;
    reg result9;

    begin
      node0_r = pixel[596];
      node0_l = ~pixel[596];
      node1_r = node0_l & pixel[263];
      node1_l = node0_l & ~pixel[263];
      node2_r = node1_l & pixel[317];
      node2_l = node1_l & ~pixel[317];
      node3_r = node2_l & pixel[326];
      node3_l = node2_l & ~pixel[326];
      node4_r = node3_l & pixel[580];
      node4_l = node3_l & ~pixel[580];
      node5_r = node4_l & pixel[466];
      node5_l = node4_l & ~pixel[466];
      node6_r = node5_l & pixel[402];
      node6_l = node5_l & ~pixel[402];
      node7_r = node6_l & pixel[234];
      node7_l = node6_l & ~pixel[234];
      node8_r = node7_l & pixel[434];
      node8_l = node7_l & ~pixel[434];
      node9_r = node8_l & pixel[544];
      node9_l = node8_l & ~pixel[544];
      node10 = node9_l;
      node11 = node9_r;
      node12_r = node8_r & pixel[522];
      node12_l = node8_r & ~pixel[522];
      node13 = node12_l;
      node14 = node12_r;
      node15_r = node7_r & pixel[375];
      node15_l = node7_r & ~pixel[375];
      node16_r = node15_l & pixel[629];
      node16_l = node15_l & ~pixel[629];
      node17 = node16_l;
      node18 = node16_r;
      node19_r = node15_r & pixel[322];
      node19_l = node15_r & ~pixel[322];
      node20 = node19_l;
      node21 = node19_r;
      node22_r = node6_r & pixel[543];
      node22_l = node6_r & ~pixel[543];
      node23_r = node22_l & pixel[245];
      node23_l = node22_l & ~pixel[245];
      node24_r = node23_l & pixel[377];
      node24_l = node23_l & ~pixel[377];
      node25 = node24_l;
      node26 = node24_r;
      node27_r = node23_r & pixel[442];
      node27_l = node23_r & ~pixel[442];
      node28 = node27_l;
      node29 = node27_r;
      node30_r = node22_r & pixel[653];
      node30_l = node22_r & ~pixel[653];
      node31_r = node30_l & pixel[406];
      node31_l = node30_l & ~pixel[406];
      node32 = node31_l;
      node33 = node31_r;
      node34_r = node30_r & pixel[400];
      node34_l = node30_r & ~pixel[400];
      node35 = node34_l;
      node36 = node34_r;
      node37_r = node5_r & pixel[513];
      node37_l = node5_r & ~pixel[513];
      node38_r = node37_l & pixel[130];
      node38_l = node37_l & ~pixel[130];
      node39_r = node38_l & pixel[515];
      node39_l = node38_l & ~pixel[515];
      node40_r = node39_l & pixel[656];
      node40_l = node39_l & ~pixel[656];
      node41 = node40_l;
      node42 = node40_r;
      node43_r = node39_r & pixel[127];
      node43_l = node39_r & ~pixel[127];
      node44 = node43_l;
      node45 = node43_r;
      node46_r = node38_r & pixel[625];
      node46_l = node38_r & ~pixel[625];
      node47_r = node46_l & pixel[297];
      node47_l = node46_l & ~pixel[297];
      node48 = node47_l;
      node49 = node47_r;
      node50_r = node46_r & pixel[457];
      node50_l = node46_r & ~pixel[457];
      node51 = node50_l;
      node52 = node50_r;
      node53_r = node37_r & pixel[403];
      node53_l = node37_r & ~pixel[403];
      node54_r = node53_l & pixel[553];
      node54_l = node53_l & ~pixel[553];
      node55_r = node54_l & pixel[347];
      node55_l = node54_l & ~pixel[347];
      node56 = node55_l;
      node57 = node55_r;
      node58_r = node54_r & pixel[551];
      node58_l = node54_r & ~pixel[551];
      node59 = node58_l;
      node60 = node58_r;
      node61_r = node53_r & pixel[601];
      node61_l = node53_r & ~pixel[601];
      node62_r = node61_l & pixel[103];
      node62_l = node61_l & ~pixel[103];
      node63 = node62_l;
      node64 = node62_r;
      node65_r = node61_r & pixel[151];
      node65_l = node61_r & ~pixel[151];
      node66 = node65_l;
      node67 = node65_r;
      node68_r = node4_r & pixel[544];
      node68_l = node4_r & ~pixel[544];
      node69_r = node68_l & pixel[321];
      node69_l = node68_l & ~pixel[321];
      node70_r = node69_l & pixel[371];
      node70_l = node69_l & ~pixel[371];
      node71_r = node70_l & pixel[496];
      node71_l = node70_l & ~pixel[496];
      node72_r = node71_l & pixel[689];
      node72_l = node71_l & ~pixel[689];
      node73 = node72_l;
      node74 = node72_r;
      node75_r = node71_r & pixel[659];
      node75_l = node71_r & ~pixel[659];
      node76 = node75_l;
      node77 = node75_r;
      node78_r = node70_r & pixel[356];
      node78_l = node70_r & ~pixel[356];
      node79_r = node78_l & pixel[376];
      node79_l = node78_l & ~pixel[376];
      node80 = node79_l;
      node81 = node79_r;
      node82_r = node78_r & pixel[599];
      node82_l = node78_r & ~pixel[599];
      node83 = node82_l;
      node84 = node82_r;
      node85_r = node69_r & pixel[568];
      node85_l = node69_r & ~pixel[568];
      node86_r = node85_l & pixel[220];
      node86_l = node85_l & ~pixel[220];
      node87_r = node86_l & pixel[485];
      node87_l = node86_l & ~pixel[485];
      node88 = node87_l;
      node89 = node87_r;
      node90 = node86_r;
      node91_r = node85_r & pixel[349];
      node91_l = node85_r & ~pixel[349];
      node92 = node91_l;
      node93_r = node91_r & pixel[411];
      node93_l = node91_r & ~pixel[411];
      node94 = node93_l;
      node95 = node93_r;
      node96_r = node68_r & pixel[322];
      node96_l = node68_r & ~pixel[322];
      node97_r = node96_l & pixel[444];
      node97_l = node96_l & ~pixel[444];
      node98_r = node97_l & pixel[370];
      node98_l = node97_l & ~pixel[370];
      node99_r = node98_l & pixel[264];
      node99_l = node98_l & ~pixel[264];
      node100 = node99_l;
      node101 = node99_r;
      node102_r = node98_r & pixel[178];
      node102_l = node98_r & ~pixel[178];
      node103 = node102_l;
      node104 = node102_r;
      node105_r = node97_r & pixel[407];
      node105_l = node97_r & ~pixel[407];
      node106_r = node105_l & pixel[436];
      node106_l = node105_l & ~pixel[436];
      node107 = node106_l;
      node108 = node106_r;
      node109 = node105_r;
      node110_r = node96_r & pixel[412];
      node110_l = node96_r & ~pixel[412];
      node111_r = node110_l & pixel[272];
      node111_l = node110_l & ~pixel[272];
      node112_r = node111_l & pixel[103];
      node112_l = node111_l & ~pixel[103];
      node113 = node112_l;
      node114 = node112_r;
      node115_r = node111_r & pixel[123];
      node115_l = node111_r & ~pixel[123];
      node116 = node115_l;
      node117 = node115_r;
      node118_r = node110_r & pixel[321];
      node118_l = node110_r & ~pixel[321];
      node119_r = node118_l & pixel[625];
      node119_l = node118_l & ~pixel[625];
      node120 = node119_l;
      node121 = node119_r;
      node122_r = node118_r & pixel[490];
      node122_l = node118_r & ~pixel[490];
      node123 = node122_l;
      node124 = node122_r;
      node125_r = node3_r & pixel[372];
      node125_l = node3_r & ~pixel[372];
      node126_r = node125_l & pixel[551];
      node126_l = node125_l & ~pixel[551];
      node127_r = node126_l & pixel[236];
      node127_l = node126_l & ~pixel[236];
      node128_r = node127_l & pixel[427];
      node128_l = node127_l & ~pixel[427];
      node129_r = node128_l & pixel[350];
      node129_l = node128_l & ~pixel[350];
      node130_r = node129_l & pixel[216];
      node130_l = node129_l & ~pixel[216];
      node131 = node130_l;
      node132 = node130_r;
      node133_r = node129_r & pixel[460];
      node133_l = node129_r & ~pixel[460];
      node134 = node133_l;
      node135 = node133_r;
      node136_r = node128_r & pixel[541];
      node136_l = node128_r & ~pixel[541];
      node137_r = node136_l & pixel[437];
      node137_l = node136_l & ~pixel[437];
      node138 = node137_l;
      node139 = node137_r;
      node140_r = node136_r & pixel[319];
      node140_l = node136_r & ~pixel[319];
      node141 = node140_l;
      node142 = node140_r;
      node143_r = node127_r & pixel[153];
      node143_l = node127_r & ~pixel[153];
      node144_r = node143_l & pixel[321];
      node144_l = node143_l & ~pixel[321];
      node145_r = node144_l & pixel[375];
      node145_l = node144_l & ~pixel[375];
      node146 = node145_l;
      node147 = node145_r;
      node148_r = node144_r & pixel[210];
      node148_l = node144_r & ~pixel[210];
      node149 = node148_l;
      node150 = node148_r;
      node151_r = node143_r & pixel[321];
      node151_l = node143_r & ~pixel[321];
      node152_r = node151_l & pixel[487];
      node152_l = node151_l & ~pixel[487];
      node153 = node152_l;
      node154 = node152_r;
      node155_r = node151_r & pixel[439];
      node155_l = node151_r & ~pixel[439];
      node156 = node155_l;
      node157 = node155_r;
      node158_r = node126_r & pixel[544];
      node158_l = node126_r & ~pixel[544];
      node159_r = node158_l & pixel[207];
      node159_l = node158_l & ~pixel[207];
      node160_r = node159_l & pixel[371];
      node160_l = node159_l & ~pixel[371];
      node161_r = node160_l & pixel[536];
      node161_l = node160_l & ~pixel[536];
      node162 = node161_l;
      node163 = node161_r;
      node164_r = node160_r & pixel[597];
      node164_l = node160_r & ~pixel[597];
      node165 = node164_l;
      node166 = node164_r;
      node167_r = node159_r & pixel[407];
      node167_l = node159_r & ~pixel[407];
      node168_r = node167_l & pixel[287];
      node168_l = node167_l & ~pixel[287];
      node169 = node168_l;
      node170 = node168_r;
      node171_r = node167_r & pixel[378];
      node171_l = node167_r & ~pixel[378];
      node172 = node171_l;
      node173 = node171_r;
      node174_r = node158_r & pixel[690];
      node174_l = node158_r & ~pixel[690];
      node175_r = node174_l & pixel[470];
      node175_l = node174_l & ~pixel[470];
      node176_r = node175_l & pixel[582];
      node176_l = node175_l & ~pixel[582];
      node177 = node176_l;
      node178 = node176_r;
      node179_r = node175_r & pixel[342];
      node179_l = node175_r & ~pixel[342];
      node180 = node179_l;
      node181 = node179_r;
      node182_r = node174_r & pixel[661];
      node182_l = node174_r & ~pixel[661];
      node183 = node182_l;
      node184_r = node182_r & pixel[152];
      node184_l = node182_r & ~pixel[152];
      node185 = node184_l;
      node186 = node184_r;
      node187_r = node125_r & pixel[207];
      node187_l = node125_r & ~pixel[207];
      node188_r = node187_l & pixel[410];
      node188_l = node187_l & ~pixel[410];
      node189_r = node188_l & pixel[402];
      node189_l = node188_l & ~pixel[402];
      node190_r = node189_l & pixel[292];
      node190_l = node189_l & ~pixel[292];
      node191_r = node190_l & pixel[213];
      node191_l = node190_l & ~pixel[213];
      node192 = node191_l;
      node193 = node191_r;
      node194_r = node190_r & pixel[602];
      node194_l = node190_r & ~pixel[602];
      node195 = node194_l;
      node196 = node194_r;
      node197_r = node189_r & pixel[274];
      node197_l = node189_r & ~pixel[274];
      node198_r = node197_l & pixel[151];
      node198_l = node197_l & ~pixel[151];
      node199 = node198_l;
      node200 = node198_r;
      node201_r = node197_r & pixel[381];
      node201_l = node197_r & ~pixel[381];
      node202 = node201_l;
      node203 = node201_r;
      node204_r = node188_r & pixel[568];
      node204_l = node188_r & ~pixel[568];
      node205_r = node204_l & pixel[93];
      node205_l = node204_l & ~pixel[93];
      node206_r = node205_l & pixel[287];
      node206_l = node205_l & ~pixel[287];
      node207 = node206_l;
      node208 = node206_r;
      node209_r = node205_r & pixel[204];
      node209_l = node205_r & ~pixel[204];
      node210 = node209_l;
      node211 = node209_r;
      node212_r = node204_r & pixel[314];
      node212_l = node204_r & ~pixel[314];
      node213_r = node212_l & pixel[327];
      node213_l = node212_l & ~pixel[327];
      node214 = node213_l;
      node215 = node213_r;
      node216_r = node212_r & pixel[547];
      node216_l = node212_r & ~pixel[547];
      node217 = node216_l;
      node218 = node216_r;
      node219_r = node187_r & pixel[343];
      node219_l = node187_r & ~pixel[343];
      node220_r = node219_l & pixel[658];
      node220_l = node219_l & ~pixel[658];
      node221_r = node220_l & pixel[519];
      node221_l = node220_l & ~pixel[519];
      node222_r = node221_l & pixel[720];
      node222_l = node221_l & ~pixel[720];
      node223 = node222_l;
      node224 = node222_r;
      node225_r = node221_r & pixel[426];
      node225_l = node221_r & ~pixel[426];
      node226 = node225_l;
      node227 = node225_r;
      node228_r = node220_r & pixel[443];
      node228_l = node220_r & ~pixel[443];
      node229 = node228_l;
      node230_r = node228_r & pixel[679];
      node230_l = node228_r & ~pixel[679];
      node231 = node230_l;
      node232 = node230_r;
      node233_r = node219_r & pixel[187];
      node233_l = node219_r & ~pixel[187];
      node234_r = node233_l & pixel[629];
      node234_l = node233_l & ~pixel[629];
      node235_r = node234_l & pixel[416];
      node235_l = node234_l & ~pixel[416];
      node236 = node235_l;
      node237 = node235_r;
      node238_r = node234_r & pixel[433];
      node238_l = node234_r & ~pixel[433];
      node239 = node238_l;
      node240 = node238_r;
      node241_r = node233_r & pixel[608];
      node241_l = node233_r & ~pixel[608];
      node242_r = node241_l & pixel[524];
      node242_l = node241_l & ~pixel[524];
      node243 = node242_l;
      node244 = node242_r;
      node245_r = node241_r & pixel[433];
      node245_l = node241_r & ~pixel[433];
      node246 = node245_l;
      node247 = node245_r;
      node248_r = node2_r & pixel[414];
      node248_l = node2_r & ~pixel[414];
      node249_r = node248_l & pixel[180];
      node249_l = node248_l & ~pixel[180];
      node250_r = node249_l & pixel[401];
      node250_l = node249_l & ~pixel[401];
      node251_r = node250_l & pixel[433];
      node251_l = node250_l & ~pixel[433];
      node252_r = node251_l & pixel[483];
      node252_l = node251_l & ~pixel[483];
      node253_r = node252_l & pixel[327];
      node253_l = node252_l & ~pixel[327];
      node254_r = node253_l & pixel[325];
      node254_l = node253_l & ~pixel[325];
      node255 = node254_l;
      node256 = node254_r;
      node257_r = node253_r & pixel[177];
      node257_l = node253_r & ~pixel[177];
      node258 = node257_l;
      node259 = node257_r;
      node260_r = node252_r & pixel[599];
      node260_l = node252_r & ~pixel[599];
      node261_r = node260_l & pixel[347];
      node261_l = node260_l & ~pixel[347];
      node262 = node261_l;
      node263 = node261_r;
      node264_r = node260_r & pixel[515];
      node264_l = node260_r & ~pixel[515];
      node265 = node264_l;
      node266 = node264_r;
      node267_r = node251_r & pixel[313];
      node267_l = node251_r & ~pixel[313];
      node268_r = node267_l & pixel[346];
      node268_l = node267_l & ~pixel[346];
      node269_r = node268_l & pixel[208];
      node269_l = node268_l & ~pixel[208];
      node270 = node269_l;
      node271 = node269_r;
      node272_r = node268_r & pixel[124];
      node272_l = node268_r & ~pixel[124];
      node273 = node272_l;
      node274 = node272_r;
      node275 = node267_r;
      node276_r = node250_r & pixel[67];
      node276_l = node250_r & ~pixel[67];
      node277_r = node276_l & pixel[293];
      node277_l = node276_l & ~pixel[293];
      node278_r = node277_l & pixel[92];
      node278_l = node277_l & ~pixel[92];
      node279_r = node278_l & pixel[597];
      node279_l = node278_l & ~pixel[597];
      node280 = node279_l;
      node281 = node279_r;
      node282 = node278_r;
      node283_r = node277_r & pixel[381];
      node283_l = node277_r & ~pixel[381];
      node284_r = node283_l & pixel[124];
      node284_l = node283_l & ~pixel[124];
      node285 = node284_l;
      node286 = node284_r;
      node287_r = node283_r & pixel[203];
      node287_l = node283_r & ~pixel[203];
      node288 = node287_l;
      node289 = node287_r;
      node290 = node276_r;
      node291_r = node249_r & pixel[497];
      node291_l = node249_r & ~pixel[497];
      node292_r = node291_l & pixel[544];
      node292_l = node291_l & ~pixel[544];
      node293_r = node292_l & pixel[156];
      node293_l = node292_l & ~pixel[156];
      node294_r = node293_l & pixel[209];
      node294_l = node293_l & ~pixel[209];
      node295_r = node294_l & pixel[273];
      node295_l = node294_l & ~pixel[273];
      node296 = node295_l;
      node297 = node295_r;
      node298_r = node294_r & pixel[653];
      node298_l = node294_r & ~pixel[653];
      node299 = node298_l;
      node300 = node298_r;
      node301_r = node293_r & pixel[467];
      node301_l = node293_r & ~pixel[467];
      node302_r = node301_l & pixel[488];
      node302_l = node301_l & ~pixel[488];
      node303 = node302_l;
      node304 = node302_r;
      node305_r = node301_r & pixel[623];
      node305_l = node301_r & ~pixel[623];
      node306 = node305_l;
      node307 = node305_r;
      node308_r = node292_r & pixel[376];
      node308_l = node292_r & ~pixel[376];
      node309_r = node308_l & pixel[301];
      node309_l = node308_l & ~pixel[301];
      node310_r = node309_l & pixel[121];
      node310_l = node309_l & ~pixel[121];
      node311 = node310_l;
      node312 = node310_r;
      node313_r = node309_r & pixel[660];
      node313_l = node309_r & ~pixel[660];
      node314 = node313_l;
      node315 = node313_r;
      node316_r = node308_r & pixel[568];
      node316_l = node308_r & ~pixel[568];
      node317_r = node316_l & pixel[341];
      node317_l = node316_l & ~pixel[341];
      node318 = node317_l;
      node319 = node317_r;
      node320_r = node316_r & pixel[495];
      node320_l = node316_r & ~pixel[495];
      node321 = node320_l;
      node322 = node320_r;
      node323_r = node291_r & pixel[325];
      node323_l = node291_r & ~pixel[325];
      node324_r = node323_l & pixel[485];
      node324_l = node323_l & ~pixel[485];
      node325_r = node324_l & pixel[185];
      node325_l = node324_l & ~pixel[185];
      node326_r = node325_l & pixel[515];
      node326_l = node325_l & ~pixel[515];
      node327 = node326_l;
      node328 = node326_r;
      node329_r = node325_r & pixel[655];
      node329_l = node325_r & ~pixel[655];
      node330 = node329_l;
      node331 = node329_r;
      node332_r = node324_r & pixel[327];
      node332_l = node324_r & ~pixel[327];
      node333_r = node332_l & pixel[660];
      node333_l = node332_l & ~pixel[660];
      node334 = node333_l;
      node335 = node333_r;
      node336_r = node332_r & pixel[212];
      node336_l = node332_r & ~pixel[212];
      node337 = node336_l;
      node338 = node336_r;
      node339_r = node323_r & pixel[265];
      node339_l = node323_r & ~pixel[265];
      node340_r = node339_l & pixel[378];
      node340_l = node339_l & ~pixel[378];
      node341_r = node340_l & pixel[429];
      node341_l = node340_l & ~pixel[429];
      node342 = node341_l;
      node343 = node341_r;
      node344_r = node340_r & pixel[406];
      node344_l = node340_r & ~pixel[406];
      node345 = node344_l;
      node346 = node344_r;
      node347_r = node339_r & pixel[378];
      node347_l = node339_r & ~pixel[378];
      node348_r = node347_l & pixel[438];
      node348_l = node347_l & ~pixel[438];
      node349 = node348_l;
      node350 = node348_r;
      node351_r = node347_r & pixel[569];
      node351_l = node347_r & ~pixel[569];
      node352 = node351_l;
      node353 = node351_r;
      node354_r = node248_r & pixel[97];
      node354_l = node248_r & ~pixel[97];
      node355_r = node354_l & pixel[121];
      node355_l = node354_l & ~pixel[121];
      node356_r = node355_l & pixel[466];
      node356_l = node355_l & ~pixel[466];
      node357_r = node356_l & pixel[518];
      node357_l = node356_l & ~pixel[518];
      node358_r = node357_l & pixel[354];
      node358_l = node357_l & ~pixel[354];
      node359_r = node358_l & pixel[541];
      node359_l = node358_l & ~pixel[541];
      node360 = node359_l;
      node361 = node359_r;
      node362_r = node358_r & pixel[239];
      node362_l = node358_r & ~pixel[239];
      node363 = node362_l;
      node364 = node362_r;
      node365_r = node357_r & pixel[185];
      node365_l = node357_r & ~pixel[185];
      node366_r = node365_l & pixel[486];
      node366_l = node365_l & ~pixel[486];
      node367 = node366_l;
      node368 = node366_r;
      node369_r = node365_r & pixel[401];
      node369_l = node365_r & ~pixel[401];
      node370 = node369_l;
      node371 = node369_r;
      node372_r = node356_r & pixel[408];
      node372_l = node356_r & ~pixel[408];
      node373_r = node372_l & pixel[348];
      node373_l = node372_l & ~pixel[348];
      node374_r = node373_l & pixel[383];
      node374_l = node373_l & ~pixel[383];
      node375 = node374_l;
      node376 = node374_r;
      node377_r = node373_r & pixel[633];
      node377_l = node373_r & ~pixel[633];
      node378 = node377_l;
      node379 = node377_r;
      node380_r = node372_r & pixel[429];
      node380_l = node372_r & ~pixel[429];
      node381_r = node380_l & pixel[456];
      node381_l = node380_l & ~pixel[456];
      node382 = node381_l;
      node383 = node381_r;
      node384_r = node380_r & pixel[153];
      node384_l = node380_r & ~pixel[153];
      node385 = node384_l;
      node386 = node384_r;
      node387_r = node355_r & pixel[660];
      node387_l = node355_r & ~pixel[660];
      node388_r = node387_l & pixel[550];
      node388_l = node387_l & ~pixel[550];
      node389_r = node388_l & pixel[445];
      node389_l = node388_l & ~pixel[445];
      node390_r = node389_l & pixel[381];
      node390_l = node389_l & ~pixel[381];
      node391 = node390_l;
      node392 = node390_r;
      node393 = node389_r;
      node394_r = node388_r & pixel[156];
      node394_l = node388_r & ~pixel[156];
      node395_r = node394_l & pixel[261];
      node395_l = node394_l & ~pixel[261];
      node396 = node395_l;
      node397 = node395_r;
      node398 = node394_r;
      node399_r = node387_r & pixel[268];
      node399_l = node387_r & ~pixel[268];
      node400_r = node399_l & pixel[293];
      node400_l = node399_l & ~pixel[293];
      node401 = node400_l;
      node402 = node400_r;
      node403_r = node399_r & pixel[469];
      node403_l = node399_r & ~pixel[469];
      node404_r = node403_l & pixel[210];
      node404_l = node403_l & ~pixel[210];
      node405 = node404_l;
      node406 = node404_r;
      node407_r = node403_r & pixel[352];
      node407_l = node403_r & ~pixel[352];
      node408 = node407_l;
      node409 = node407_r;
      node410 = node354_r;
      node411_r = node1_r & pixel[432];
      node411_l = node1_r & ~pixel[432];
      node412_r = node411_l & pixel[181];
      node412_l = node411_l & ~pixel[181];
      node413_r = node412_l & pixel[483];
      node413_l = node412_l & ~pixel[483];
      node414_r = node413_l & pixel[404];
      node414_l = node413_l & ~pixel[404];
      node415_r = node414_l & pixel[430];
      node415_l = node414_l & ~pixel[430];
      node416_r = node415_l & pixel[152];
      node416_l = node415_l & ~pixel[152];
      node417_r = node416_l & pixel[542];
      node417_l = node416_l & ~pixel[542];
      node418_r = node417_l & pixel[350];
      node418_l = node417_l & ~pixel[350];
      node419 = node418_l;
      node420 = node418_r;
      node421_r = node417_r & pixel[241];
      node421_l = node417_r & ~pixel[241];
      node422 = node421_l;
      node423 = node421_r;
      node424_r = node416_r & pixel[523];
      node424_l = node416_r & ~pixel[523];
      node425_r = node424_l & pixel[127];
      node425_l = node424_l & ~pixel[127];
      node426 = node425_l;
      node427 = node425_r;
      node428_r = node424_r & pixel[321];
      node428_l = node424_r & ~pixel[321];
      node429 = node428_l;
      node430 = node428_r;
      node431_r = node415_r & pixel[68];
      node431_l = node415_r & ~pixel[68];
      node432_r = node431_l & pixel[461];
      node432_l = node431_l & ~pixel[461];
      node433_r = node432_l & pixel[385];
      node433_l = node432_l & ~pixel[385];
      node434 = node433_l;
      node435 = node433_r;
      node436_r = node432_r & pixel[440];
      node436_l = node432_r & ~pixel[440];
      node437 = node436_l;
      node438 = node436_r;
      node439 = node431_r;
      node440_r = node414_r & pixel[523];
      node440_l = node414_r & ~pixel[523];
      node441_r = node440_l & pixel[178];
      node441_l = node440_l & ~pixel[178];
      node442_r = node441_l & pixel[632];
      node442_l = node441_l & ~pixel[632];
      node443_r = node442_l & pixel[212];
      node443_l = node442_l & ~pixel[212];
      node444 = node443_l;
      node445 = node443_r;
      node446_r = node442_r & pixel[324];
      node446_l = node442_r & ~pixel[324];
      node447 = node446_l;
      node448 = node446_r;
      node449_r = node441_r & pixel[486];
      node449_l = node441_r & ~pixel[486];
      node450_r = node449_l & pixel[374];
      node450_l = node449_l & ~pixel[374];
      node451 = node450_l;
      node452 = node450_r;
      node453_r = node449_r & pixel[185];
      node453_l = node449_r & ~pixel[185];
      node454 = node453_l;
      node455 = node453_r;
      node456_r = node440_r & pixel[286];
      node456_l = node440_r & ~pixel[286];
      node457_r = node456_l & pixel[102];
      node457_l = node456_l & ~pixel[102];
      node458_r = node457_l & pixel[201];
      node458_l = node457_l & ~pixel[201];
      node459 = node458_l;
      node460 = node458_r;
      node461 = node457_r;
      node462_r = node456_r & pixel[409];
      node462_l = node456_r & ~pixel[409];
      node463_r = node462_l & pixel[211];
      node463_l = node462_l & ~pixel[211];
      node464 = node463_l;
      node465 = node463_r;
      node466_r = node462_r & pixel[400];
      node466_l = node462_r & ~pixel[400];
      node467 = node466_l;
      node468 = node466_r;
      node469_r = node413_r & pixel[331];
      node469_l = node413_r & ~pixel[331];
      node470_r = node469_l & pixel[569];
      node470_l = node469_l & ~pixel[569];
      node471_r = node470_l & pixel[491];
      node471_l = node470_l & ~pixel[491];
      node472_r = node471_l & pixel[486];
      node472_l = node471_l & ~pixel[486];
      node473_r = node472_l & pixel[380];
      node473_l = node472_l & ~pixel[380];
      node474 = node473_l;
      node475 = node473_r;
      node476_r = node472_r & pixel[205];
      node476_l = node472_r & ~pixel[205];
      node477 = node476_l;
      node478 = node476_r;
      node479_r = node471_r & pixel[747];
      node479_l = node471_r & ~pixel[747];
      node480_r = node479_l & pixel[159];
      node480_l = node479_l & ~pixel[159];
      node481 = node480_l;
      node482 = node480_r;
      node483 = node479_r;
      node484_r = node470_r & pixel[130];
      node484_l = node470_r & ~pixel[130];
      node485_r = node484_l & pixel[463];
      node485_l = node484_l & ~pixel[463];
      node486_r = node485_l & pixel[177];
      node486_l = node485_l & ~pixel[177];
      node487 = node486_l;
      node488 = node486_r;
      node489_r = node485_r & pixel[599];
      node489_l = node485_r & ~pixel[599];
      node490 = node489_l;
      node491 = node489_r;
      node492_r = node484_r & pixel[320];
      node492_l = node484_r & ~pixel[320];
      node493 = node492_l;
      node494_r = node492_r & pixel[412];
      node494_l = node492_r & ~pixel[412];
      node495 = node494_l;
      node496 = node494_r;
      node497_r = node469_r & pixel[381];
      node497_l = node469_r & ~pixel[381];
      node498_r = node497_l & pixel[121];
      node498_l = node497_l & ~pixel[121];
      node499_r = node498_l & pixel[526];
      node499_l = node498_l & ~pixel[526];
      node500_r = node499_l & pixel[573];
      node500_l = node499_l & ~pixel[573];
      node501 = node500_l;
      node502 = node500_r;
      node503_r = node499_r & pixel[314];
      node503_l = node499_r & ~pixel[314];
      node504 = node503_l;
      node505 = node503_r;
      node506 = node498_r;
      node507_r = node497_r & pixel[513];
      node507_l = node497_r & ~pixel[513];
      node508_r = node507_l & pixel[188];
      node508_l = node507_l & ~pixel[188];
      node509 = node508_l;
      node510 = node508_r;
      node511_r = node507_r & pixel[179];
      node511_l = node507_r & ~pixel[179];
      node512_r = node511_l & pixel[269];
      node512_l = node511_l & ~pixel[269];
      node513 = node512_l;
      node514 = node512_r;
      node515_r = node511_r & pixel[215];
      node515_l = node511_r & ~pixel[215];
      node516 = node515_l;
      node517 = node515_r;
      node518_r = node412_r & pixel[212];
      node518_l = node412_r & ~pixel[212];
      node519_r = node518_l & pixel[515];
      node519_l = node518_l & ~pixel[515];
      node520_r = node519_l & pixel[631];
      node520_l = node519_l & ~pixel[631];
      node521_r = node520_l & pixel[268];
      node521_l = node520_l & ~pixel[268];
      node522_r = node521_l & pixel[541];
      node522_l = node521_l & ~pixel[541];
      node523_r = node522_l & pixel[402];
      node523_l = node522_l & ~pixel[402];
      node524 = node523_l;
      node525 = node523_r;
      node526_r = node522_r & pixel[660];
      node526_l = node522_r & ~pixel[660];
      node527 = node526_l;
      node528 = node526_r;
      node529_r = node521_r & pixel[717];
      node529_l = node521_r & ~pixel[717];
      node530_r = node529_l & pixel[578];
      node530_l = node529_l & ~pixel[578];
      node531 = node530_l;
      node532 = node530_r;
      node533 = node529_r;
      node534_r = node520_r & pixel[495];
      node534_l = node520_r & ~pixel[495];
      node535_r = node534_l & pixel[547];
      node535_l = node534_l & ~pixel[547];
      node536_r = node535_l & pixel[520];
      node536_l = node535_l & ~pixel[520];
      node537 = node536_l;
      node538 = node536_r;
      node539_r = node535_r & pixel[353];
      node539_l = node535_r & ~pixel[353];
      node540 = node539_l;
      node541 = node539_r;
      node542_r = node534_r & pixel[456];
      node542_l = node534_r & ~pixel[456];
      node543_r = node542_l & pixel[157];
      node543_l = node542_l & ~pixel[157];
      node544 = node543_l;
      node545 = node543_r;
      node546_r = node542_r & pixel[434];
      node546_l = node542_r & ~pixel[434];
      node547 = node546_l;
      node548 = node546_r;
      node549_r = node519_r & pixel[186];
      node549_l = node519_r & ~pixel[186];
      node550_r = node549_l & pixel[656];
      node550_l = node549_l & ~pixel[656];
      node551_r = node550_l & pixel[272];
      node551_l = node550_l & ~pixel[272];
      node552_r = node551_l & pixel[121];
      node552_l = node551_l & ~pixel[121];
      node553 = node552_l;
      node554 = node552_r;
      node555_r = node551_r & pixel[100];
      node555_l = node551_r & ~pixel[100];
      node556 = node555_l;
      node557 = node555_r;
      node558_r = node550_r & pixel[322];
      node558_l = node550_r & ~pixel[322];
      node559_r = node558_l & pixel[518];
      node559_l = node558_l & ~pixel[518];
      node560 = node559_l;
      node561 = node559_r;
      node562_r = node558_r & pixel[384];
      node562_l = node558_r & ~pixel[384];
      node563 = node562_l;
      node564 = node562_r;
      node565_r = node549_r & pixel[407];
      node565_l = node549_r & ~pixel[407];
      node566_r = node565_l & pixel[328];
      node566_l = node565_l & ~pixel[328];
      node567_r = node566_l & pixel[569];
      node567_l = node566_l & ~pixel[569];
      node568 = node567_l;
      node569 = node567_r;
      node570_r = node566_r & pixel[125];
      node570_l = node566_r & ~pixel[125];
      node571 = node570_l;
      node572 = node570_r;
      node573_r = node565_r & pixel[403];
      node573_l = node565_r & ~pixel[403];
      node574_r = node573_l & pixel[433];
      node574_l = node573_l & ~pixel[433];
      node575 = node574_l;
      node576 = node574_r;
      node577_r = node573_r & pixel[655];
      node577_l = node573_r & ~pixel[655];
      node578 = node577_l;
      node579 = node577_r;
      node580_r = node518_r & pixel[155];
      node580_l = node518_r & ~pixel[155];
      node581_r = node580_l & pixel[428];
      node581_l = node580_l & ~pixel[428];
      node582_r = node581_l & pixel[298];
      node582_l = node581_l & ~pixel[298];
      node583_r = node582_l & pixel[188];
      node583_l = node582_l & ~pixel[188];
      node584_r = node583_l & pixel[491];
      node584_l = node583_l & ~pixel[491];
      node585 = node584_l;
      node586 = node584_r;
      node587_r = node583_r & pixel[488];
      node587_l = node583_r & ~pixel[488];
      node588 = node587_l;
      node589 = node587_r;
      node590_r = node582_r & pixel[430];
      node590_l = node582_r & ~pixel[430];
      node591_r = node590_l & pixel[349];
      node591_l = node590_l & ~pixel[349];
      node592 = node591_l;
      node593 = node591_r;
      node594_r = node590_r & pixel[570];
      node594_l = node590_r & ~pixel[570];
      node595 = node594_l;
      node596 = node594_r;
      node597_r = node581_r & pixel[598];
      node597_l = node581_r & ~pixel[598];
      node598_r = node597_l & pixel[653];
      node598_l = node597_l & ~pixel[653];
      node599_r = node598_l & pixel[487];
      node599_l = node598_l & ~pixel[487];
      node600 = node599_l;
      node601 = node599_r;
      node602_r = node598_r & pixel[435];
      node602_l = node598_r & ~pixel[435];
      node603 = node602_l;
      node604 = node602_r;
      node605_r = node597_r & pixel[376];
      node605_l = node597_r & ~pixel[376];
      node606_r = node605_l & pixel[485];
      node606_l = node605_l & ~pixel[485];
      node607 = node606_l;
      node608 = node606_r;
      node609_r = node605_r & pixel[546];
      node609_l = node605_r & ~pixel[546];
      node610 = node609_l;
      node611 = node609_r;
      node612_r = node580_r & pixel[463];
      node612_l = node580_r & ~pixel[463];
      node613_r = node612_l & pixel[569];
      node613_l = node612_l & ~pixel[569];
      node614_r = node613_l & pixel[356];
      node614_l = node613_l & ~pixel[356];
      node615_r = node614_l & pixel[331];
      node615_l = node614_l & ~pixel[331];
      node616 = node615_l;
      node617 = node615_r;
      node618_r = node614_r & pixel[542];
      node618_l = node614_r & ~pixel[542];
      node619 = node618_l;
      node620 = node618_r;
      node621_r = node613_r & pixel[322];
      node621_l = node613_r & ~pixel[322];
      node622_r = node621_l & pixel[350];
      node622_l = node621_l & ~pixel[350];
      node623 = node622_l;
      node624 = node622_r;
      node625_r = node621_r & pixel[350];
      node625_l = node621_r & ~pixel[350];
      node626 = node625_l;
      node627 = node625_r;
      node628_r = node612_r & pixel[296];
      node628_l = node612_r & ~pixel[296];
      node629_r = node628_l & pixel[101];
      node629_l = node628_l & ~pixel[101];
      node630_r = node629_l & pixel[406];
      node630_l = node629_l & ~pixel[406];
      node631 = node630_l;
      node632 = node630_r;
      node633_r = node629_r & pixel[378];
      node633_l = node629_r & ~pixel[378];
      node634 = node633_l;
      node635 = node633_r;
      node636_r = node628_r & pixel[351];
      node636_l = node628_r & ~pixel[351];
      node637_r = node636_l & pixel[571];
      node637_l = node636_l & ~pixel[571];
      node638 = node637_l;
      node639 = node637_r;
      node640_r = node636_r & pixel[625];
      node640_l = node636_r & ~pixel[625];
      node641 = node640_l;
      node642 = node640_r;
      node643_r = node411_r & pixel[127];
      node643_l = node411_r & ~pixel[127];
      node644_r = node643_l & pixel[183];
      node644_l = node643_l & ~pixel[183];
      node645_r = node644_l & pixel[294];
      node645_l = node644_l & ~pixel[294];
      node646_r = node645_l & pixel[162];
      node646_l = node645_l & ~pixel[162];
      node647_r = node646_l & pixel[212];
      node647_l = node646_l & ~pixel[212];
      node648_r = node647_l & pixel[551];
      node648_l = node647_l & ~pixel[551];
      node649_r = node648_l & pixel[267];
      node649_l = node648_l & ~pixel[267];
      node650 = node649_l;
      node651 = node649_r;
      node652_r = node648_r & pixel[572];
      node652_l = node648_r & ~pixel[572];
      node653 = node652_l;
      node654 = node652_r;
      node655_r = node647_r & pixel[209];
      node655_l = node647_r & ~pixel[209];
      node656_r = node655_l & pixel[323];
      node656_l = node655_l & ~pixel[323];
      node657 = node656_l;
      node658 = node656_r;
      node659_r = node655_r & pixel[409];
      node659_l = node655_r & ~pixel[409];
      node660 = node659_l;
      node661 = node659_r;
      node662_r = node646_r & pixel[409];
      node662_l = node646_r & ~pixel[409];
      node663_r = node662_l & pixel[244];
      node663_l = node662_l & ~pixel[244];
      node664 = node663_l;
      node665_r = node663_r & pixel[427];
      node665_l = node663_r & ~pixel[427];
      node666 = node665_l;
      node667 = node665_r;
      node668_r = node662_r & pixel[622];
      node668_l = node662_r & ~pixel[622];
      node669_r = node668_l & pixel[428];
      node669_l = node668_l & ~pixel[428];
      node670 = node669_l;
      node671 = node669_r;
      node672 = node668_r;
      node673_r = node645_r & pixel[526];
      node673_l = node645_r & ~pixel[526];
      node674_r = node673_l & pixel[345];
      node674_l = node673_l & ~pixel[345];
      node675_r = node674_l & pixel[290];
      node675_l = node674_l & ~pixel[290];
      node676_r = node675_l & pixel[325];
      node676_l = node675_l & ~pixel[325];
      node677 = node676_l;
      node678 = node676_r;
      node679_r = node675_r & pixel[343];
      node679_l = node675_r & ~pixel[343];
      node680 = node679_l;
      node681 = node679_r;
      node682_r = node674_r & pixel[239];
      node682_l = node674_r & ~pixel[239];
      node683_r = node682_l & pixel[382];
      node683_l = node682_l & ~pixel[382];
      node684 = node683_l;
      node685 = node683_r;
      node686_r = node682_r & pixel[352];
      node686_l = node682_r & ~pixel[352];
      node687 = node686_l;
      node688 = node686_r;
      node689_r = node673_r & pixel[632];
      node689_l = node673_r & ~pixel[632];
      node690_r = node689_l & pixel[662];
      node690_l = node689_l & ~pixel[662];
      node691_r = node690_l & pixel[299];
      node691_l = node690_l & ~pixel[299];
      node692 = node691_l;
      node693 = node691_r;
      node694_r = node690_r & pixel[609];
      node694_l = node690_r & ~pixel[609];
      node695 = node694_l;
      node696 = node694_r;
      node697_r = node689_r & pixel[543];
      node697_l = node689_r & ~pixel[543];
      node698_r = node697_l & pixel[515];
      node698_l = node697_l & ~pixel[515];
      node699 = node698_l;
      node700 = node698_r;
      node701_r = node697_r & pixel[435];
      node701_l = node697_r & ~pixel[435];
      node702 = node701_l;
      node703 = node701_r;
      node704_r = node644_r & pixel[158];
      node704_l = node644_r & ~pixel[158];
      node705_r = node704_l & pixel[409];
      node705_l = node704_l & ~pixel[409];
      node706_r = node705_l & pixel[219];
      node706_l = node705_l & ~pixel[219];
      node707_r = node706_l & pixel[380];
      node707_l = node706_l & ~pixel[380];
      node708_r = node707_l & pixel[324];
      node708_l = node707_l & ~pixel[324];
      node709 = node708_l;
      node710 = node708_r;
      node711_r = node707_r & pixel[599];
      node711_l = node707_r & ~pixel[599];
      node712 = node711_l;
      node713 = node711_r;
      node714_r = node706_r & pixel[570];
      node714_l = node706_r & ~pixel[570];
      node715_r = node714_l & pixel[298];
      node715_l = node714_l & ~pixel[298];
      node716 = node715_l;
      node717 = node715_r;
      node718_r = node714_r & pixel[343];
      node718_l = node714_r & ~pixel[343];
      node719 = node718_l;
      node720 = node718_r;
      node721_r = node705_r & pixel[441];
      node721_l = node705_r & ~pixel[441];
      node722_r = node721_l & pixel[372];
      node722_l = node721_l & ~pixel[372];
      node723_r = node722_l & pixel[155];
      node723_l = node722_l & ~pixel[155];
      node724 = node723_l;
      node725 = node723_r;
      node726_r = node722_r & pixel[219];
      node726_l = node722_r & ~pixel[219];
      node727 = node726_l;
      node728 = node726_r;
      node729_r = node721_r & pixel[518];
      node729_l = node721_r & ~pixel[518];
      node730_r = node729_l & pixel[397];
      node730_l = node729_l & ~pixel[397];
      node731 = node730_l;
      node732 = node730_r;
      node733_r = node729_r & pixel[268];
      node733_l = node729_r & ~pixel[268];
      node734 = node733_l;
      node735 = node733_r;
      node736_r = node704_r & pixel[652];
      node736_l = node704_r & ~pixel[652];
      node737_r = node736_l & pixel[484];
      node737_l = node736_l & ~pixel[484];
      node738_r = node737_l & pixel[518];
      node738_l = node737_l & ~pixel[518];
      node739_r = node738_l & pixel[571];
      node739_l = node738_l & ~pixel[571];
      node740 = node739_l;
      node741 = node739_r;
      node742_r = node738_r & pixel[405];
      node742_l = node738_r & ~pixel[405];
      node743 = node742_l;
      node744 = node742_r;
      node745_r = node737_r & pixel[686];
      node745_l = node737_r & ~pixel[686];
      node746_r = node745_l & pixel[609];
      node746_l = node745_l & ~pixel[609];
      node747 = node746_l;
      node748 = node746_r;
      node749_r = node745_r & pixel[607];
      node749_l = node745_r & ~pixel[607];
      node750 = node749_l;
      node751 = node749_r;
      node752_r = node736_r & pixel[512];
      node752_l = node736_r & ~pixel[512];
      node753_r = node752_l & pixel[325];
      node753_l = node752_l & ~pixel[325];
      node754_r = node753_l & pixel[298];
      node754_l = node753_l & ~pixel[298];
      node755 = node754_l;
      node756 = node754_r;
      node757_r = node753_r & pixel[597];
      node757_l = node753_r & ~pixel[597];
      node758 = node757_l;
      node759 = node757_r;
      node760_r = node752_r & pixel[497];
      node760_l = node752_r & ~pixel[497];
      node761_r = node760_l & pixel[352];
      node761_l = node760_l & ~pixel[352];
      node762 = node761_l;
      node763 = node761_r;
      node764_r = node760_r & pixel[357];
      node764_l = node760_r & ~pixel[357];
      node765 = node764_l;
      node766 = node764_r;
      node767_r = node643_r & pixel[269];
      node767_l = node643_r & ~pixel[269];
      node768_r = node767_l & pixel[486];
      node768_l = node767_l & ~pixel[486];
      node769_r = node768_l & pixel[103];
      node769_l = node768_l & ~pixel[103];
      node770_r = node769_l & pixel[628];
      node770_l = node769_l & ~pixel[628];
      node771_r = node770_l & pixel[99];
      node771_l = node770_l & ~pixel[99];
      node772_r = node771_l & pixel[540];
      node772_l = node771_l & ~pixel[540];
      node773 = node772_l;
      node774 = node772_r;
      node775_r = node771_r & pixel[494];
      node775_l = node771_r & ~pixel[494];
      node776 = node775_l;
      node777 = node775_r;
      node778_r = node770_r & pixel[460];
      node778_l = node770_r & ~pixel[460];
      node779_r = node778_l & pixel[329];
      node779_l = node778_l & ~pixel[329];
      node780 = node779_l;
      node781 = node779_r;
      node782_r = node778_r & pixel[296];
      node782_l = node778_r & ~pixel[296];
      node783 = node782_l;
      node784 = node782_r;
      node785 = node769_r;
      node786_r = node768_r & pixel[655];
      node786_l = node768_r & ~pixel[655];
      node787_r = node786_l & pixel[271];
      node787_l = node786_l & ~pixel[271];
      node788_r = node787_l & pixel[656];
      node788_l = node787_l & ~pixel[656];
      node789_r = node788_l & pixel[543];
      node789_l = node788_l & ~pixel[543];
      node790 = node789_l;
      node791 = node789_r;
      node792_r = node788_r & pixel[409];
      node792_l = node788_r & ~pixel[409];
      node793 = node792_l;
      node794 = node792_r;
      node795_r = node787_r & pixel[456];
      node795_l = node787_r & ~pixel[456];
      node796_r = node795_l & pixel[550];
      node796_l = node795_l & ~pixel[550];
      node797 = node796_l;
      node798 = node796_r;
      node799_r = node795_r & pixel[600];
      node799_l = node795_r & ~pixel[600];
      node800 = node799_l;
      node801 = node799_r;
      node802_r = node786_r & pixel[659];
      node802_l = node786_r & ~pixel[659];
      node803_r = node802_l & pixel[214];
      node803_l = node802_l & ~pixel[214];
      node804_r = node803_l & pixel[184];
      node804_l = node803_l & ~pixel[184];
      node805 = node804_l;
      node806 = node804_r;
      node807_r = node803_r & pixel[461];
      node807_l = node803_r & ~pixel[461];
      node808 = node807_l;
      node809 = node807_r;
      node810_r = node802_r & pixel[230];
      node810_l = node802_r & ~pixel[230];
      node811_r = node810_l & pixel[238];
      node811_l = node810_l & ~pixel[238];
      node812 = node811_l;
      node813 = node811_r;
      node814 = node810_r;
      node815_r = node767_r & pixel[356];
      node815_l = node767_r & ~pixel[356];
      node816_r = node815_l & pixel[481];
      node816_l = node815_l & ~pixel[481];
      node817_r = node816_l & pixel[484];
      node817_l = node816_l & ~pixel[484];
      node818_r = node817_l & pixel[583];
      node818_l = node817_l & ~pixel[583];
      node819_r = node818_l & pixel[434];
      node819_l = node818_l & ~pixel[434];
      node820 = node819_l;
      node821 = node819_r;
      node822 = node818_r;
      node823_r = node817_r & pixel[399];
      node823_l = node817_r & ~pixel[399];
      node824_r = node823_l & pixel[519];
      node824_l = node823_l & ~pixel[519];
      node825 = node824_l;
      node826 = node824_r;
      node827_r = node823_r & pixel[547];
      node827_l = node823_r & ~pixel[547];
      node828 = node827_l;
      node829 = node827_r;
      node830_r = node816_r & pixel[566];
      node830_l = node816_r & ~pixel[566];
      node831_r = node830_l & pixel[592];
      node831_l = node830_l & ~pixel[592];
      node832 = node831_l;
      node833 = node831_r;
      node834 = node830_r;
      node835_r = node815_r & pixel[433];
      node835_l = node815_r & ~pixel[433];
      node836_r = node835_l & pixel[185];
      node836_l = node835_l & ~pixel[185];
      node837_r = node836_l & pixel[607];
      node837_l = node836_l & ~pixel[607];
      node838 = node837_l;
      node839_r = node837_r & pixel[100];
      node839_l = node837_r & ~pixel[100];
      node840 = node839_l;
      node841 = node839_r;
      node842_r = node836_r & pixel[178];
      node842_l = node836_r & ~pixel[178];
      node843 = node842_l;
      node844_r = node842_r & pixel[491];
      node844_l = node842_r & ~pixel[491];
      node845 = node844_l;
      node846 = node844_r;
      node847_r = node835_r & pixel[572];
      node847_l = node835_r & ~pixel[572];
      node848_r = node847_l & pixel[344];
      node848_l = node847_l & ~pixel[344];
      node849 = node848_l;
      node850_r = node848_r & pixel[152];
      node850_l = node848_r & ~pixel[152];
      node851 = node850_l;
      node852 = node850_r;
      node853_r = node847_r & pixel[213];
      node853_l = node847_r & ~pixel[213];
      node854 = node853_l;
      node855_r = node853_r & pixel[347];
      node855_l = node853_r & ~pixel[347];
      node856 = node855_l;
      node857 = node855_r;
      node858_r = node0_r & pixel[352];
      node858_l = node0_r & ~pixel[352];
      node859_r = node858_l & pixel[316];
      node859_l = node858_l & ~pixel[316];
      node860_r = node859_l & pixel[318];
      node860_l = node859_l & ~pixel[318];
      node861_r = node860_l & pixel[517];
      node861_l = node860_l & ~pixel[517];
      node862_r = node861_l & pixel[151];
      node862_l = node861_l & ~pixel[151];
      node863_r = node862_l & pixel[484];
      node863_l = node862_l & ~pixel[484];
      node864_r = node863_l & pixel[292];
      node864_l = node863_l & ~pixel[292];
      node865_r = node864_l & pixel[378];
      node865_l = node864_l & ~pixel[378];
      node866_r = node865_l & pixel[499];
      node866_l = node865_l & ~pixel[499];
      node867 = node866_l;
      node868 = node866_r;
      node869_r = node865_r & pixel[515];
      node869_l = node865_r & ~pixel[515];
      node870 = node869_l;
      node871 = node869_r;
      node872_r = node864_r & pixel[385];
      node872_l = node864_r & ~pixel[385];
      node873_r = node872_l & pixel[201];
      node873_l = node872_l & ~pixel[201];
      node874 = node873_l;
      node875 = node873_r;
      node876_r = node872_r & pixel[434];
      node876_l = node872_r & ~pixel[434];
      node877 = node876_l;
      node878 = node876_r;
      node879_r = node863_r & pixel[347];
      node879_l = node863_r & ~pixel[347];
      node880_r = node879_l & pixel[579];
      node880_l = node879_l & ~pixel[579];
      node881_r = node880_l & pixel[342];
      node881_l = node880_l & ~pixel[342];
      node882 = node881_l;
      node883 = node881_r;
      node884_r = node880_r & pixel[548];
      node884_l = node880_r & ~pixel[548];
      node885 = node884_l;
      node886 = node884_r;
      node887_r = node879_r & pixel[436];
      node887_l = node879_r & ~pixel[436];
      node888_r = node887_l & pixel[329];
      node888_l = node887_l & ~pixel[329];
      node889 = node888_l;
      node890 = node888_r;
      node891_r = node887_r & pixel[327];
      node891_l = node887_r & ~pixel[327];
      node892 = node891_l;
      node893 = node891_r;
      node894_r = node862_r & pixel[658];
      node894_l = node862_r & ~pixel[658];
      node895_r = node894_l & pixel[397];
      node895_l = node894_l & ~pixel[397];
      node896_r = node895_l & pixel[539];
      node896_l = node895_l & ~pixel[539];
      node897_r = node896_l & pixel[322];
      node897_l = node896_l & ~pixel[322];
      node898 = node897_l;
      node899 = node897_r;
      node900_r = node896_r & pixel[490];
      node900_l = node896_r & ~pixel[490];
      node901 = node900_l;
      node902 = node900_r;
      node903_r = node895_r & pixel[594];
      node903_l = node895_r & ~pixel[594];
      node904_r = node903_l & pixel[623];
      node904_l = node903_l & ~pixel[623];
      node905 = node904_l;
      node906 = node904_r;
      node907 = node903_r;
      node908_r = node894_r & pixel[349];
      node908_l = node894_r & ~pixel[349];
      node909_r = node908_l & pixel[342];
      node909_l = node908_l & ~pixel[342];
      node910_r = node909_l & pixel[265];
      node910_l = node909_l & ~pixel[265];
      node911 = node910_l;
      node912 = node910_r;
      node913_r = node909_r & pixel[436];
      node913_l = node909_r & ~pixel[436];
      node914 = node913_l;
      node915 = node913_r;
      node916_r = node908_r & pixel[357];
      node916_l = node908_r & ~pixel[357];
      node917_r = node916_l & pixel[294];
      node917_l = node916_l & ~pixel[294];
      node918 = node917_l;
      node919 = node917_r;
      node920_r = node916_r & pixel[437];
      node920_l = node916_r & ~pixel[437];
      node921 = node920_l;
      node922 = node920_r;
      node923_r = node861_r & pixel[322];
      node923_l = node861_r & ~pixel[322];
      node924_r = node923_l & pixel[706];
      node924_l = node923_l & ~pixel[706];
      node925_r = node924_l & pixel[655];
      node925_l = node924_l & ~pixel[655];
      node926_r = node925_l & pixel[164];
      node926_l = node925_l & ~pixel[164];
      node927_r = node926_l & pixel[127];
      node927_l = node926_l & ~pixel[127];
      node928 = node927_l;
      node929 = node927_r;
      node930_r = node926_r & pixel[427];
      node930_l = node926_r & ~pixel[427];
      node931 = node930_l;
      node932 = node930_r;
      node933_r = node925_r & pixel[495];
      node933_l = node925_r & ~pixel[495];
      node934_r = node933_l & pixel[432];
      node934_l = node933_l & ~pixel[432];
      node935 = node934_l;
      node936 = node934_r;
      node937_r = node933_r & pixel[528];
      node937_l = node933_r & ~pixel[528];
      node938 = node937_l;
      node939 = node937_r;
      node940_r = node924_r & pixel[348];
      node940_l = node924_r & ~pixel[348];
      node941 = node940_l;
      node942 = node940_r;
      node943_r = node923_r & pixel[132];
      node943_l = node923_r & ~pixel[132];
      node944_r = node943_l & pixel[384];
      node944_l = node943_l & ~pixel[384];
      node945_r = node944_l & pixel[128];
      node945_l = node944_l & ~pixel[128];
      node946_r = node945_l & pixel[180];
      node946_l = node945_l & ~pixel[180];
      node947 = node946_l;
      node948 = node946_r;
      node949_r = node945_r & pixel[179];
      node949_l = node945_r & ~pixel[179];
      node950 = node949_l;
      node951 = node949_r;
      node952_r = node944_r & pixel[409];
      node952_l = node944_r & ~pixel[409];
      node953_r = node952_l & pixel[216];
      node953_l = node952_l & ~pixel[216];
      node954 = node953_l;
      node955 = node953_r;
      node956_r = node952_r & pixel[428];
      node956_l = node952_r & ~pixel[428];
      node957 = node956_l;
      node958 = node956_r;
      node959_r = node943_r & pixel[622];
      node959_l = node943_r & ~pixel[622];
      node960_r = node959_l & pixel[459];
      node960_l = node959_l & ~pixel[459];
      node961_r = node960_l & pixel[457];
      node961_l = node960_l & ~pixel[457];
      node962 = node961_l;
      node963 = node961_r;
      node964_r = node960_r & pixel[426];
      node964_l = node960_r & ~pixel[426];
      node965 = node964_l;
      node966 = node964_r;
      node967_r = node959_r & pixel[402];
      node967_l = node959_r & ~pixel[402];
      node968_r = node967_l & pixel[217];
      node968_l = node967_l & ~pixel[217];
      node969 = node968_l;
      node970 = node968_r;
      node971_r = node967_r & pixel[578];
      node971_l = node967_r & ~pixel[578];
      node972 = node971_l;
      node973 = node971_r;
      node974_r = node860_r & pixel[484];
      node974_l = node860_r & ~pixel[484];
      node975_r = node974_l & pixel[543];
      node975_l = node974_l & ~pixel[543];
      node976_r = node975_l & pixel[357];
      node976_l = node975_l & ~pixel[357];
      node977_r = node976_l & pixel[122];
      node977_l = node976_l & ~pixel[122];
      node978_r = node977_l & pixel[178];
      node978_l = node977_l & ~pixel[178];
      node979_r = node978_l & pixel[414];
      node979_l = node978_l & ~pixel[414];
      node980 = node979_l;
      node981 = node979_r;
      node982_r = node978_r & pixel[175];
      node982_l = node978_r & ~pixel[175];
      node983 = node982_l;
      node984 = node982_r;
      node985_r = node977_r & pixel[296];
      node985_l = node977_r & ~pixel[296];
      node986_r = node985_l & pixel[176];
      node986_l = node985_l & ~pixel[176];
      node987 = node986_l;
      node988 = node986_r;
      node989 = node985_r;
      node990_r = node976_r & pixel[486];
      node990_l = node976_r & ~pixel[486];
      node991_r = node990_l & pixel[147];
      node991_l = node990_l & ~pixel[147];
      node992_r = node991_l & pixel[292];
      node992_l = node991_l & ~pixel[292];
      node993 = node992_l;
      node994 = node992_r;
      node995 = node991_r;
      node996_r = node990_r & pixel[456];
      node996_l = node990_r & ~pixel[456];
      node997_r = node996_l & pixel[377];
      node997_l = node996_l & ~pixel[377];
      node998 = node997_l;
      node999 = node997_r;
      node1000 = node996_r;
      node1001_r = node975_r & pixel[509];
      node1001_l = node975_r & ~pixel[509];
      node1002_r = node1001_l & pixel[354];
      node1002_l = node1001_l & ~pixel[354];
      node1003_r = node1002_l & pixel[157];
      node1003_l = node1002_l & ~pixel[157];
      node1004_r = node1003_l & pixel[358];
      node1004_l = node1003_l & ~pixel[358];
      node1005 = node1004_l;
      node1006 = node1004_r;
      node1007_r = node1003_r & pixel[383];
      node1007_l = node1003_r & ~pixel[383];
      node1008 = node1007_l;
      node1009 = node1007_r;
      node1010_r = node1002_r & pixel[656];
      node1010_l = node1002_r & ~pixel[656];
      node1011_r = node1010_l & pixel[432];
      node1011_l = node1010_l & ~pixel[432];
      node1012 = node1011_l;
      node1013 = node1011_r;
      node1014_r = node1010_r & pixel[495];
      node1014_l = node1010_r & ~pixel[495];
      node1015 = node1014_l;
      node1016 = node1014_r;
      node1017_r = node1001_r & pixel[344];
      node1017_l = node1001_r & ~pixel[344];
      node1018_r = node1017_l & pixel[441];
      node1018_l = node1017_l & ~pixel[441];
      node1019_r = node1018_l & pixel[384];
      node1019_l = node1018_l & ~pixel[384];
      node1020 = node1019_l;
      node1021 = node1019_r;
      node1022_r = node1018_r & pixel[623];
      node1022_l = node1018_r & ~pixel[623];
      node1023 = node1022_l;
      node1024 = node1022_r;
      node1025_r = node1017_r & pixel[432];
      node1025_l = node1017_r & ~pixel[432];
      node1026_r = node1025_l & pixel[462];
      node1026_l = node1025_l & ~pixel[462];
      node1027 = node1026_l;
      node1028 = node1026_r;
      node1029_r = node1025_r & pixel[565];
      node1029_l = node1025_r & ~pixel[565];
      node1030 = node1029_l;
      node1031 = node1029_r;
      node1032_r = node974_r & pixel[461];
      node1032_l = node974_r & ~pixel[461];
      node1033_r = node1032_l & pixel[243];
      node1033_l = node1032_l & ~pixel[243];
      node1034_r = node1033_l & pixel[655];
      node1034_l = node1033_l & ~pixel[655];
      node1035_r = node1034_l & pixel[273];
      node1035_l = node1034_l & ~pixel[273];
      node1036_r = node1035_l & pixel[245];
      node1036_l = node1035_l & ~pixel[245];
      node1037 = node1036_l;
      node1038 = node1036_r;
      node1039_r = node1035_r & pixel[374];
      node1039_l = node1035_r & ~pixel[374];
      node1040 = node1039_l;
      node1041 = node1039_r;
      node1042_r = node1034_r & pixel[374];
      node1042_l = node1034_r & ~pixel[374];
      node1043_r = node1042_l & pixel[357];
      node1043_l = node1042_l & ~pixel[357];
      node1044 = node1043_l;
      node1045 = node1043_r;
      node1046_r = node1042_r & pixel[379];
      node1046_l = node1042_r & ~pixel[379];
      node1047 = node1046_l;
      node1048 = node1046_r;
      node1049_r = node1033_r & pixel[405];
      node1049_l = node1033_r & ~pixel[405];
      node1050_r = node1049_l & pixel[384];
      node1050_l = node1049_l & ~pixel[384];
      node1051_r = node1050_l & pixel[191];
      node1051_l = node1050_l & ~pixel[191];
      node1052 = node1051_l;
      node1053 = node1051_r;
      node1054_r = node1050_r & pixel[428];
      node1054_l = node1050_r & ~pixel[428];
      node1055 = node1054_l;
      node1056 = node1054_r;
      node1057_r = node1049_r & pixel[220];
      node1057_l = node1049_r & ~pixel[220];
      node1058_r = node1057_l & pixel[429];
      node1058_l = node1057_l & ~pixel[429];
      node1059 = node1058_l;
      node1060 = node1058_r;
      node1061_r = node1057_r & pixel[359];
      node1061_l = node1057_r & ~pixel[359];
      node1062 = node1061_l;
      node1063 = node1061_r;
      node1064_r = node1032_r & pixel[467];
      node1064_l = node1032_r & ~pixel[467];
      node1065_r = node1064_l & pixel[207];
      node1065_l = node1064_l & ~pixel[207];
      node1066_r = node1065_l & pixel[157];
      node1066_l = node1065_l & ~pixel[157];
      node1067_r = node1066_l & pixel[331];
      node1067_l = node1066_l & ~pixel[331];
      node1068 = node1067_l;
      node1069 = node1067_r;
      node1070_r = node1066_r & pixel[244];
      node1070_l = node1066_r & ~pixel[244];
      node1071 = node1070_l;
      node1072 = node1070_r;
      node1073_r = node1065_r & pixel[541];
      node1073_l = node1065_r & ~pixel[541];
      node1074_r = node1073_l & pixel[345];
      node1074_l = node1073_l & ~pixel[345];
      node1075 = node1074_l;
      node1076 = node1074_r;
      node1077_r = node1073_r & pixel[348];
      node1077_l = node1073_r & ~pixel[348];
      node1078 = node1077_l;
      node1079 = node1077_r;
      node1080_r = node1064_r & pixel[622];
      node1080_l = node1064_r & ~pixel[622];
      node1081_r = node1080_l & pixel[299];
      node1081_l = node1080_l & ~pixel[299];
      node1082_r = node1081_l & pixel[216];
      node1082_l = node1081_l & ~pixel[216];
      node1083 = node1082_l;
      node1084 = node1082_r;
      node1085_r = node1081_r & pixel[629];
      node1085_l = node1081_r & ~pixel[629];
      node1086 = node1085_l;
      node1087 = node1085_r;
      node1088_r = node1080_r & pixel[128];
      node1088_l = node1080_r & ~pixel[128];
      node1089_r = node1088_l & pixel[578];
      node1089_l = node1088_l & ~pixel[578];
      node1090 = node1089_l;
      node1091 = node1089_r;
      node1092_r = node1088_r & pixel[131];
      node1092_l = node1088_r & ~pixel[131];
      node1093 = node1092_l;
      node1094 = node1092_r;
      node1095_r = node859_r & pixel[425];
      node1095_l = node859_r & ~pixel[425];
      node1096_r = node1095_l & pixel[469];
      node1096_l = node1095_l & ~pixel[469];
      node1097_r = node1096_l & pixel[330];
      node1097_l = node1096_l & ~pixel[330];
      node1098_r = node1097_l & pixel[353];
      node1098_l = node1097_l & ~pixel[353];
      node1099_r = node1098_l & pixel[383];
      node1099_l = node1098_l & ~pixel[383];
      node1100_r = node1099_l & pixel[126];
      node1100_l = node1099_l & ~pixel[126];
      node1101_r = node1100_l & pixel[471];
      node1101_l = node1100_l & ~pixel[471];
      node1102 = node1101_l;
      node1103 = node1101_r;
      node1104_r = node1100_r & pixel[130];
      node1104_l = node1100_r & ~pixel[130];
      node1105 = node1104_l;
      node1106 = node1104_r;
      node1107_r = node1099_r & pixel[372];
      node1107_l = node1099_r & ~pixel[372];
      node1108_r = node1107_l & pixel[275];
      node1108_l = node1107_l & ~pixel[275];
      node1109 = node1108_l;
      node1110 = node1108_r;
      node1111_r = node1107_r & pixel[553];
      node1111_l = node1107_r & ~pixel[553];
      node1112 = node1111_l;
      node1113 = node1111_r;
      node1114_r = node1098_r & pixel[467];
      node1114_l = node1098_r & ~pixel[467];
      node1115_r = node1114_l & pixel[567];
      node1115_l = node1114_l & ~pixel[567];
      node1116_r = node1115_l & pixel[185];
      node1116_l = node1115_l & ~pixel[185];
      node1117 = node1116_l;
      node1118 = node1116_r;
      node1119_r = node1115_r & pixel[357];
      node1119_l = node1115_r & ~pixel[357];
      node1120 = node1119_l;
      node1121 = node1119_r;
      node1122_r = node1114_r & pixel[344];
      node1122_l = node1114_r & ~pixel[344];
      node1123_r = node1122_l & pixel[681];
      node1123_l = node1122_l & ~pixel[681];
      node1124 = node1123_l;
      node1125 = node1123_r;
      node1126_r = node1122_r & pixel[434];
      node1126_l = node1122_r & ~pixel[434];
      node1127 = node1126_l;
      node1128 = node1126_r;
      node1129_r = node1097_r & pixel[382];
      node1129_l = node1097_r & ~pixel[382];
      node1130_r = node1129_l & pixel[491];
      node1130_l = node1129_l & ~pixel[491];
      node1131_r = node1130_l & pixel[455];
      node1131_l = node1130_l & ~pixel[455];
      node1132_r = node1131_l & pixel[548];
      node1132_l = node1131_l & ~pixel[548];
      node1133 = node1132_l;
      node1134 = node1132_r;
      node1135_r = node1131_r & pixel[162];
      node1135_l = node1131_r & ~pixel[162];
      node1136 = node1135_l;
      node1137 = node1135_r;
      node1138_r = node1130_r & pixel[277];
      node1138_l = node1130_r & ~pixel[277];
      node1139_r = node1138_l & pixel[270];
      node1139_l = node1138_l & ~pixel[270];
      node1140 = node1139_l;
      node1141 = node1139_r;
      node1142_r = node1138_r & pixel[521];
      node1142_l = node1138_r & ~pixel[521];
      node1143 = node1142_l;
      node1144 = node1142_r;
      node1145_r = node1129_r & pixel[706];
      node1145_l = node1129_r & ~pixel[706];
      node1146_r = node1145_l & pixel[399];
      node1146_l = node1145_l & ~pixel[399];
      node1147_r = node1146_l & pixel[373];
      node1147_l = node1146_l & ~pixel[373];
      node1148 = node1147_l;
      node1149 = node1147_r;
      node1150_r = node1146_r & pixel[516];
      node1150_l = node1146_r & ~pixel[516];
      node1151 = node1150_l;
      node1152 = node1150_r;
      node1153_r = node1145_r & pixel[487];
      node1153_l = node1145_r & ~pixel[487];
      node1154_r = node1153_l & pixel[405];
      node1154_l = node1153_l & ~pixel[405];
      node1155 = node1154_l;
      node1156 = node1154_r;
      node1157_r = node1153_r & pixel[657];
      node1157_l = node1153_r & ~pixel[657];
      node1158 = node1157_l;
      node1159 = node1157_r;
      node1160_r = node1096_r & pixel[463];
      node1160_l = node1096_r & ~pixel[463];
      node1161_r = node1160_l & pixel[407];
      node1161_l = node1160_l & ~pixel[407];
      node1162_r = node1161_l & pixel[145];
      node1162_l = node1161_l & ~pixel[145];
      node1163_r = node1162_l & pixel[507];
      node1163_l = node1162_l & ~pixel[507];
      node1164_r = node1163_l & pixel[648];
      node1164_l = node1163_l & ~pixel[648];
      node1165 = node1164_l;
      node1166 = node1164_r;
      node1167 = node1163_r;
      node1168 = node1162_r;
      node1169_r = node1161_r & pixel[328];
      node1169_l = node1161_r & ~pixel[328];
      node1170_r = node1169_l & pixel[99];
      node1170_l = node1169_l & ~pixel[99];
      node1171_r = node1170_l & pixel[105];
      node1171_l = node1170_l & ~pixel[105];
      node1172 = node1171_l;
      node1173 = node1171_r;
      node1174_r = node1170_r & pixel[624];
      node1174_l = node1170_r & ~pixel[624];
      node1175 = node1174_l;
      node1176 = node1174_r;
      node1177_r = node1169_r & pixel[321];
      node1177_l = node1169_r & ~pixel[321];
      node1178_r = node1177_l & pixel[623];
      node1178_l = node1177_l & ~pixel[623];
      node1179 = node1178_l;
      node1180 = node1178_r;
      node1181 = node1177_r;
      node1182_r = node1160_r & pixel[655];
      node1182_l = node1160_r & ~pixel[655];
      node1183_r = node1182_l & pixel[213];
      node1183_l = node1182_l & ~pixel[213];
      node1184_r = node1183_l & pixel[259];
      node1184_l = node1183_l & ~pixel[259];
      node1185_r = node1184_l & pixel[70];
      node1185_l = node1184_l & ~pixel[70];
      node1186 = node1185_l;
      node1187 = node1185_r;
      node1188_r = node1184_r & pixel[356];
      node1188_l = node1184_r & ~pixel[356];
      node1189 = node1188_l;
      node1190 = node1188_r;
      node1191_r = node1183_r & pixel[320];
      node1191_l = node1183_r & ~pixel[320];
      node1192_r = node1191_l & pixel[358];
      node1192_l = node1191_l & ~pixel[358];
      node1193 = node1192_l;
      node1194 = node1192_r;
      node1195_r = node1191_r & pixel[400];
      node1195_l = node1191_r & ~pixel[400];
      node1196 = node1195_l;
      node1197 = node1195_r;
      node1198_r = node1182_r & pixel[600];
      node1198_l = node1182_r & ~pixel[600];
      node1199_r = node1198_l & pixel[357];
      node1199_l = node1198_l & ~pixel[357];
      node1200_r = node1199_l & pixel[516];
      node1200_l = node1199_l & ~pixel[516];
      node1201 = node1200_l;
      node1202 = node1200_r;
      node1203 = node1199_r;
      node1204_r = node1198_r & pixel[526];
      node1204_l = node1198_r & ~pixel[526];
      node1205_r = node1204_l & pixel[158];
      node1205_l = node1204_l & ~pixel[158];
      node1206 = node1205_l;
      node1207 = node1205_r;
      node1208_r = node1204_r & pixel[606];
      node1208_l = node1204_r & ~pixel[606];
      node1209 = node1208_l;
      node1210 = node1208_r;
      node1211_r = node1095_r & pixel[462];
      node1211_l = node1095_r & ~pixel[462];
      node1212_r = node1211_l & pixel[73];
      node1212_l = node1211_l & ~pixel[73];
      node1213_r = node1212_l & pixel[70];
      node1213_l = node1212_l & ~pixel[70];
      node1214_r = node1213_l & pixel[381];
      node1214_l = node1213_l & ~pixel[381];
      node1215_r = node1214_l & pixel[693];
      node1215_l = node1214_l & ~pixel[693];
      node1216_r = node1215_l & pixel[243];
      node1216_l = node1215_l & ~pixel[243];
      node1217 = node1216_l;
      node1218 = node1216_r;
      node1219_r = node1215_r & pixel[690];
      node1219_l = node1215_r & ~pixel[690];
      node1220 = node1219_l;
      node1221 = node1219_r;
      node1222_r = node1214_r & pixel[407];
      node1222_l = node1214_r & ~pixel[407];
      node1223_r = node1222_l & pixel[629];
      node1223_l = node1222_l & ~pixel[629];
      node1224 = node1223_l;
      node1225 = node1223_r;
      node1226_r = node1222_r & pixel[383];
      node1226_l = node1222_r & ~pixel[383];
      node1227 = node1226_l;
      node1228 = node1226_r;
      node1229 = node1213_r;
      node1230 = node1212_r;
      node1231_r = node1211_r & pixel[378];
      node1231_l = node1211_r & ~pixel[378];
      node1232_r = node1231_l & pixel[300];
      node1232_l = node1231_l & ~pixel[300];
      node1233_r = node1232_l & pixel[689];
      node1233_l = node1232_l & ~pixel[689];
      node1234_r = node1233_l & pixel[368];
      node1234_l = node1233_l & ~pixel[368];
      node1235 = node1234_l;
      node1236 = node1234_r;
      node1237 = node1233_r;
      node1238_r = node1232_r & pixel[268];
      node1238_l = node1232_r & ~pixel[268];
      node1239_r = node1238_l & pixel[246];
      node1239_l = node1238_l & ~pixel[246];
      node1240_r = node1239_l & pixel[511];
      node1240_l = node1239_l & ~pixel[511];
      node1241 = node1240_l;
      node1242 = node1240_r;
      node1243_r = node1239_r & pixel[128];
      node1243_l = node1239_r & ~pixel[128];
      node1244 = node1243_l;
      node1245 = node1243_r;
      node1246_r = node1238_r & pixel[472];
      node1246_l = node1238_r & ~pixel[472];
      node1247_r = node1246_l & pixel[375];
      node1247_l = node1246_l & ~pixel[375];
      node1248 = node1247_l;
      node1249 = node1247_r;
      node1250 = node1246_r;
      node1251_r = node1231_r & pixel[631];
      node1251_l = node1231_r & ~pixel[631];
      node1252_r = node1251_l & pixel[693];
      node1252_l = node1251_l & ~pixel[693];
      node1253 = node1252_l;
      node1254 = node1252_r;
      node1255_r = node1251_r & pixel[608];
      node1255_l = node1251_r & ~pixel[608];
      node1256_r = node1255_l & pixel[373];
      node1256_l = node1255_l & ~pixel[373];
      node1257 = node1256_l;
      node1258 = node1256_r;
      node1259_r = node1255_r & pixel[301];
      node1259_l = node1255_r & ~pixel[301];
      node1260 = node1259_l;
      node1261 = node1259_r;
      node1262_r = node858_r & pixel[376];
      node1262_l = node858_r & ~pixel[376];
      node1263_r = node1262_l & pixel[124];
      node1263_l = node1262_l & ~pixel[124];
      node1264_r = node1263_l & pixel[235];
      node1264_l = node1263_l & ~pixel[235];
      node1265_r = node1264_l & pixel[154];
      node1265_l = node1264_l & ~pixel[154];
      node1266_r = node1265_l & pixel[320];
      node1266_l = node1265_l & ~pixel[320];
      node1267_r = node1266_l & pixel[265];
      node1267_l = node1266_l & ~pixel[265];
      node1268_r = node1267_l & pixel[374];
      node1268_l = node1267_l & ~pixel[374];
      node1269_r = node1268_l & pixel[546];
      node1269_l = node1268_l & ~pixel[546];
      node1270 = node1269_l;
      node1271 = node1269_r;
      node1272_r = node1268_r & pixel[510];
      node1272_l = node1268_r & ~pixel[510];
      node1273 = node1272_l;
      node1274 = node1272_r;
      node1275_r = node1267_r & pixel[484];
      node1275_l = node1267_r & ~pixel[484];
      node1276_r = node1275_l & pixel[522];
      node1276_l = node1275_l & ~pixel[522];
      node1277 = node1276_l;
      node1278 = node1276_r;
      node1279_r = node1275_r & pixel[626];
      node1279_l = node1275_r & ~pixel[626];
      node1280 = node1279_l;
      node1281 = node1279_r;
      node1282_r = node1266_r & pixel[372];
      node1282_l = node1266_r & ~pixel[372];
      node1283_r = node1282_l & pixel[290];
      node1283_l = node1282_l & ~pixel[290];
      node1284_r = node1283_l & pixel[524];
      node1284_l = node1283_l & ~pixel[524];
      node1285 = node1284_l;
      node1286 = node1284_r;
      node1287_r = node1283_r & pixel[350];
      node1287_l = node1283_r & ~pixel[350];
      node1288 = node1287_l;
      node1289 = node1287_r;
      node1290_r = node1282_r & pixel[130];
      node1290_l = node1282_r & ~pixel[130];
      node1291_r = node1290_l & pixel[262];
      node1291_l = node1290_l & ~pixel[262];
      node1292 = node1291_l;
      node1293 = node1291_r;
      node1294_r = node1290_r & pixel[269];
      node1294_l = node1290_r & ~pixel[269];
      node1295 = node1294_l;
      node1296 = node1294_r;
      node1297_r = node1265_r & pixel[348];
      node1297_l = node1265_r & ~pixel[348];
      node1298_r = node1297_l & pixel[569];
      node1298_l = node1297_l & ~pixel[569];
      node1299_r = node1298_l & pixel[438];
      node1299_l = node1298_l & ~pixel[438];
      node1300_r = node1299_l & pixel[150];
      node1300_l = node1299_l & ~pixel[150];
      node1301 = node1300_l;
      node1302 = node1300_r;
      node1303_r = node1299_r & pixel[403];
      node1303_l = node1299_r & ~pixel[403];
      node1304 = node1303_l;
      node1305 = node1303_r;
      node1306_r = node1298_r & pixel[349];
      node1306_l = node1298_r & ~pixel[349];
      node1307_r = node1306_l & pixel[321];
      node1307_l = node1306_l & ~pixel[321];
      node1308 = node1307_l;
      node1309 = node1307_r;
      node1310_r = node1306_r & pixel[460];
      node1310_l = node1306_r & ~pixel[460];
      node1311 = node1310_l;
      node1312 = node1310_r;
      node1313_r = node1297_r & pixel[433];
      node1313_l = node1297_r & ~pixel[433];
      node1314_r = node1313_l & pixel[289];
      node1314_l = node1313_l & ~pixel[289];
      node1315_r = node1314_l & pixel[237];
      node1315_l = node1314_l & ~pixel[237];
      node1316 = node1315_l;
      node1317 = node1315_r;
      node1318_r = node1314_r & pixel[466];
      node1318_l = node1314_r & ~pixel[466];
      node1319 = node1318_l;
      node1320 = node1318_r;
      node1321_r = node1313_r & pixel[456];
      node1321_l = node1313_r & ~pixel[456];
      node1322_r = node1321_l & pixel[651];
      node1322_l = node1321_l & ~pixel[651];
      node1323 = node1322_l;
      node1324 = node1322_r;
      node1325 = node1321_r;
      node1326_r = node1264_r & pixel[544];
      node1326_l = node1264_r & ~pixel[544];
      node1327_r = node1326_l & pixel[435];
      node1327_l = node1326_l & ~pixel[435];
      node1328_r = node1327_l & pixel[388];
      node1328_l = node1327_l & ~pixel[388];
      node1329_r = node1328_l & pixel[455];
      node1329_l = node1328_l & ~pixel[455];
      node1330_r = node1329_l & pixel[272];
      node1330_l = node1329_l & ~pixel[272];
      node1331 = node1330_l;
      node1332 = node1330_r;
      node1333_r = node1329_r & pixel[271];
      node1333_l = node1329_r & ~pixel[271];
      node1334 = node1333_l;
      node1335 = node1333_r;
      node1336 = node1328_r;
      node1337_r = node1327_r & pixel[232];
      node1337_l = node1327_r & ~pixel[232];
      node1338_r = node1337_l & pixel[537];
      node1338_l = node1337_l & ~pixel[537];
      node1339_r = node1338_l & pixel[540];
      node1339_l = node1338_l & ~pixel[540];
      node1340 = node1339_l;
      node1341 = node1339_r;
      node1342_r = node1338_r & pixel[525];
      node1342_l = node1338_r & ~pixel[525];
      node1343 = node1342_l;
      node1344 = node1342_r;
      node1345_r = node1337_r & pixel[438];
      node1345_l = node1337_r & ~pixel[438];
      node1346_r = node1345_l & pixel[513];
      node1346_l = node1345_l & ~pixel[513];
      node1347 = node1346_l;
      node1348 = node1346_r;
      node1349_r = node1345_r & pixel[495];
      node1349_l = node1345_r & ~pixel[495];
      node1350 = node1349_l;
      node1351 = node1349_r;
      node1352_r = node1326_r & pixel[709];
      node1352_l = node1326_r & ~pixel[709];
      node1353_r = node1352_l & pixel[413];
      node1353_l = node1352_l & ~pixel[413];
      node1354_r = node1353_l & pixel[274];
      node1354_l = node1353_l & ~pixel[274];
      node1355_r = node1354_l & pixel[163];
      node1355_l = node1354_l & ~pixel[163];
      node1356 = node1355_l;
      node1357 = node1355_r;
      node1358_r = node1354_r & pixel[511];
      node1358_l = node1354_r & ~pixel[511];
      node1359 = node1358_l;
      node1360 = node1358_r;
      node1361_r = node1353_r & pixel[517];
      node1361_l = node1353_r & ~pixel[517];
      node1362_r = node1361_l & pixel[370];
      node1362_l = node1361_l & ~pixel[370];
      node1363 = node1362_l;
      node1364 = node1362_r;
      node1365_r = node1361_r & pixel[241];
      node1365_l = node1361_r & ~pixel[241];
      node1366 = node1365_l;
      node1367 = node1365_r;
      node1368_r = node1352_r & pixel[490];
      node1368_l = node1352_r & ~pixel[490];
      node1369_r = node1368_l & pixel[320];
      node1369_l = node1368_l & ~pixel[320];
      node1370 = node1369_l;
      node1371 = node1369_r;
      node1372_r = node1368_r & pixel[456];
      node1372_l = node1368_r & ~pixel[456];
      node1373_r = node1372_l & pixel[621];
      node1373_l = node1372_l & ~pixel[621];
      node1374 = node1373_l;
      node1375 = node1373_r;
      node1376_r = node1372_r & pixel[329];
      node1376_l = node1372_r & ~pixel[329];
      node1377 = node1376_l;
      node1378 = node1376_r;
      node1379_r = node1263_r & pixel[349];
      node1379_l = node1263_r & ~pixel[349];
      node1380_r = node1379_l & pixel[330];
      node1380_l = node1379_l & ~pixel[330];
      node1381_r = node1380_l & pixel[384];
      node1381_l = node1380_l & ~pixel[384];
      node1382_r = node1381_l & pixel[264];
      node1382_l = node1381_l & ~pixel[264];
      node1383_r = node1382_l & pixel[568];
      node1383_l = node1382_l & ~pixel[568];
      node1384_r = node1383_l & pixel[120];
      node1384_l = node1383_l & ~pixel[120];
      node1385 = node1384_l;
      node1386 = node1384_r;
      node1387_r = node1383_r & pixel[246];
      node1387_l = node1383_r & ~pixel[246];
      node1388 = node1387_l;
      node1389 = node1387_r;
      node1390_r = node1382_r & pixel[490];
      node1390_l = node1382_r & ~pixel[490];
      node1391_r = node1390_l & pixel[237];
      node1391_l = node1390_l & ~pixel[237];
      node1392 = node1391_l;
      node1393 = node1391_r;
      node1394_r = node1390_r & pixel[246];
      node1394_l = node1390_r & ~pixel[246];
      node1395 = node1394_l;
      node1396 = node1394_r;
      node1397_r = node1381_r & pixel[434];
      node1397_l = node1381_r & ~pixel[434];
      node1398_r = node1397_l & pixel[373];
      node1398_l = node1397_l & ~pixel[373];
      node1399_r = node1398_l & pixel[323];
      node1399_l = node1398_l & ~pixel[323];
      node1400 = node1399_l;
      node1401 = node1399_r;
      node1402 = node1398_r;
      node1403_r = node1397_r & pixel[488];
      node1403_l = node1397_r & ~pixel[488];
      node1404_r = node1403_l & pixel[122];
      node1404_l = node1403_l & ~pixel[122];
      node1405 = node1404_l;
      node1406 = node1404_r;
      node1407_r = node1403_r & pixel[327];
      node1407_l = node1403_r & ~pixel[327];
      node1408 = node1407_l;
      node1409 = node1407_r;
      node1410_r = node1380_r & pixel[608];
      node1410_l = node1380_r & ~pixel[608];
      node1411_r = node1410_l & pixel[621];
      node1411_l = node1410_l & ~pixel[621];
      node1412_r = node1411_l & pixel[317];
      node1412_l = node1411_l & ~pixel[317];
      node1413_r = node1412_l & pixel[549];
      node1413_l = node1412_l & ~pixel[549];
      node1414 = node1413_l;
      node1415 = node1413_r;
      node1416_r = node1412_r & pixel[158];
      node1416_l = node1412_r & ~pixel[158];
      node1417 = node1416_l;
      node1418 = node1416_r;
      node1419 = node1411_r;
      node1420_r = node1410_r & pixel[401];
      node1420_l = node1410_r & ~pixel[401];
      node1421 = node1420_l;
      node1422 = node1420_r;
      node1423_r = node1379_r & pixel[490];
      node1423_l = node1379_r & ~pixel[490];
      node1424_r = node1423_l & pixel[516];
      node1424_l = node1423_l & ~pixel[516];
      node1425_r = node1424_l & pixel[296];
      node1425_l = node1424_l & ~pixel[296];
      node1426_r = node1425_l & pixel[260];
      node1426_l = node1425_l & ~pixel[260];
      node1427_r = node1426_l & pixel[464];
      node1427_l = node1426_l & ~pixel[464];
      node1428 = node1427_l;
      node1429 = node1427_r;
      node1430_r = node1426_r & pixel[271];
      node1430_l = node1426_r & ~pixel[271];
      node1431 = node1430_l;
      node1432 = node1430_r;
      node1433_r = node1425_r & pixel[541];
      node1433_l = node1425_r & ~pixel[541];
      node1434_r = node1433_l & pixel[443];
      node1434_l = node1433_l & ~pixel[443];
      node1435 = node1434_l;
      node1436 = node1434_r;
      node1437_r = node1433_r & pixel[298];
      node1437_l = node1433_r & ~pixel[298];
      node1438 = node1437_l;
      node1439 = node1437_r;
      node1440_r = node1424_r & pixel[405];
      node1440_l = node1424_r & ~pixel[405];
      node1441_r = node1440_l & pixel[636];
      node1441_l = node1440_l & ~pixel[636];
      node1442_r = node1441_l & pixel[538];
      node1442_l = node1441_l & ~pixel[538];
      node1443 = node1442_l;
      node1444 = node1442_r;
      node1445 = node1441_r;
      node1446_r = node1440_r & pixel[292];
      node1446_l = node1440_r & ~pixel[292];
      node1447_r = node1446_l & pixel[262];
      node1447_l = node1446_l & ~pixel[262];
      node1448 = node1447_l;
      node1449 = node1447_r;
      node1450_r = node1446_r & pixel[212];
      node1450_l = node1446_r & ~pixel[212];
      node1451 = node1450_l;
      node1452 = node1450_r;
      node1453_r = node1423_r & pixel[553];
      node1453_l = node1423_r & ~pixel[553];
      node1454_r = node1453_l & pixel[296];
      node1454_l = node1453_l & ~pixel[296];
      node1455_r = node1454_l & pixel[496];
      node1455_l = node1454_l & ~pixel[496];
      node1456 = node1455_l;
      node1457 = node1455_r;
      node1458_r = node1454_r & pixel[602];
      node1458_l = node1454_r & ~pixel[602];
      node1459 = node1458_l;
      node1460_r = node1458_r & pixel[469];
      node1460_l = node1458_r & ~pixel[469];
      node1461 = node1460_l;
      node1462 = node1460_r;
      node1463 = node1453_r;
      node1464_r = node1262_r & pixel[180];
      node1464_l = node1262_r & ~pixel[180];
      node1465_r = node1464_l & pixel[460];
      node1465_l = node1464_l & ~pixel[460];
      node1466_r = node1465_l & pixel[265];
      node1466_l = node1465_l & ~pixel[265];
      node1467_r = node1466_l & pixel[324];
      node1467_l = node1466_l & ~pixel[324];
      node1468_r = node1467_l & pixel[453];
      node1468_l = node1467_l & ~pixel[453];
      node1469_r = node1468_l & pixel[357];
      node1469_l = node1468_l & ~pixel[357];
      node1470_r = node1469_l & pixel[125];
      node1470_l = node1469_l & ~pixel[125];
      node1471 = node1470_l;
      node1472 = node1470_r;
      node1473_r = node1469_r & pixel[469];
      node1473_l = node1469_r & ~pixel[469];
      node1474 = node1473_l;
      node1475 = node1473_r;
      node1476 = node1468_r;
      node1477_r = node1467_r & pixel[626];
      node1477_l = node1467_r & ~pixel[626];
      node1478_r = node1477_l & pixel[127];
      node1478_l = node1477_l & ~pixel[127];
      node1479_r = node1478_l & pixel[380];
      node1479_l = node1478_l & ~pixel[380];
      node1480 = node1479_l;
      node1481 = node1479_r;
      node1482_r = node1478_r & pixel[599];
      node1482_l = node1478_r & ~pixel[599];
      node1483 = node1482_l;
      node1484 = node1482_r;
      node1485_r = node1477_r & pixel[303];
      node1485_l = node1477_r & ~pixel[303];
      node1486_r = node1485_l & pixel[555];
      node1486_l = node1485_l & ~pixel[555];
      node1487 = node1486_l;
      node1488 = node1486_r;
      node1489_r = node1485_r & pixel[189];
      node1489_l = node1485_r & ~pixel[189];
      node1490 = node1489_l;
      node1491 = node1489_r;
      node1492_r = node1466_r & pixel[488];
      node1492_l = node1466_r & ~pixel[488];
      node1493_r = node1492_l & pixel[326];
      node1493_l = node1492_l & ~pixel[326];
      node1494_r = node1493_l & pixel[122];
      node1494_l = node1493_l & ~pixel[122];
      node1495_r = node1494_l & pixel[219];
      node1495_l = node1494_l & ~pixel[219];
      node1496 = node1495_l;
      node1497 = node1495_r;
      node1498 = node1494_r;
      node1499_r = node1493_r & pixel[331];
      node1499_l = node1493_r & ~pixel[331];
      node1500_r = node1499_l & pixel[485];
      node1500_l = node1499_l & ~pixel[485];
      node1501 = node1500_l;
      node1502 = node1500_r;
      node1503_r = node1499_r & pixel[539];
      node1503_l = node1499_r & ~pixel[539];
      node1504 = node1503_l;
      node1505 = node1503_r;
      node1506_r = node1492_r & pixel[512];
      node1506_l = node1492_r & ~pixel[512];
      node1507_r = node1506_l & pixel[630];
      node1507_l = node1506_l & ~pixel[630];
      node1508_r = node1507_l & pixel[461];
      node1508_l = node1507_l & ~pixel[461];
      node1509 = node1508_l;
      node1510 = node1508_r;
      node1511 = node1507_r;
      node1512_r = node1506_r & pixel[348];
      node1512_l = node1506_r & ~pixel[348];
      node1513 = node1512_l;
      node1514_r = node1512_r & pixel[358];
      node1514_l = node1512_r & ~pixel[358];
      node1515 = node1514_l;
      node1516 = node1514_r;
      node1517_r = node1465_r & pixel[320];
      node1517_l = node1465_r & ~pixel[320];
      node1518_r = node1517_l & pixel[237];
      node1518_l = node1517_l & ~pixel[237];
      node1519_r = node1518_l & pixel[551];
      node1519_l = node1518_l & ~pixel[551];
      node1520_r = node1519_l & pixel[322];
      node1520_l = node1519_l & ~pixel[322];
      node1521_r = node1520_l & pixel[217];
      node1521_l = node1520_l & ~pixel[217];
      node1522 = node1521_l;
      node1523 = node1521_r;
      node1524_r = node1520_r & pixel[406];
      node1524_l = node1520_r & ~pixel[406];
      node1525 = node1524_l;
      node1526 = node1524_r;
      node1527_r = node1519_r & pixel[470];
      node1527_l = node1519_r & ~pixel[470];
      node1528_r = node1527_l & pixel[570];
      node1528_l = node1527_l & ~pixel[570];
      node1529 = node1528_l;
      node1530 = node1528_r;
      node1531_r = node1527_r & pixel[299];
      node1531_l = node1527_r & ~pixel[299];
      node1532 = node1531_l;
      node1533 = node1531_r;
      node1534_r = node1518_r & pixel[536];
      node1534_l = node1518_r & ~pixel[536];
      node1535_r = node1534_l & pixel[410];
      node1535_l = node1534_l & ~pixel[410];
      node1536_r = node1535_l & pixel[567];
      node1536_l = node1535_l & ~pixel[567];
      node1537 = node1536_l;
      node1538 = node1536_r;
      node1539_r = node1535_r & pixel[291];
      node1539_l = node1535_r & ~pixel[291];
      node1540 = node1539_l;
      node1541 = node1539_r;
      node1542_r = node1534_r & pixel[512];
      node1542_l = node1534_r & ~pixel[512];
      node1543 = node1542_l;
      node1544 = node1542_r;
      node1545_r = node1517_r & pixel[271];
      node1545_l = node1517_r & ~pixel[271];
      node1546_r = node1545_l & pixel[411];
      node1546_l = node1545_l & ~pixel[411];
      node1547_r = node1546_l & pixel[326];
      node1547_l = node1546_l & ~pixel[326];
      node1548_r = node1547_l & pixel[269];
      node1548_l = node1547_l & ~pixel[269];
      node1549 = node1548_l;
      node1550 = node1548_r;
      node1551_r = node1547_r & pixel[152];
      node1551_l = node1547_r & ~pixel[152];
      node1552 = node1551_l;
      node1553 = node1551_r;
      node1554_r = node1546_r & pixel[273];
      node1554_l = node1546_r & ~pixel[273];
      node1555_r = node1554_l & pixel[217];
      node1555_l = node1554_l & ~pixel[217];
      node1556 = node1555_l;
      node1557 = node1555_r;
      node1558_r = node1554_r & pixel[574];
      node1558_l = node1554_r & ~pixel[574];
      node1559 = node1558_l;
      node1560 = node1558_r;
      node1561_r = node1545_r & pixel[374];
      node1561_l = node1545_r & ~pixel[374];
      node1562_r = node1561_l & pixel[407];
      node1562_l = node1561_l & ~pixel[407];
      node1563_r = node1562_l & pixel[193];
      node1563_l = node1562_l & ~pixel[193];
      node1564 = node1563_l;
      node1565 = node1563_r;
      node1566_r = node1562_r & pixel[292];
      node1566_l = node1562_r & ~pixel[292];
      node1567 = node1566_l;
      node1568 = node1566_r;
      node1569_r = node1561_r & pixel[214];
      node1569_l = node1561_r & ~pixel[214];
      node1570_r = node1569_l & pixel[410];
      node1570_l = node1569_l & ~pixel[410];
      node1571 = node1570_l;
      node1572 = node1570_r;
      node1573_r = node1569_r & pixel[210];
      node1573_l = node1569_r & ~pixel[210];
      node1574 = node1573_l;
      node1575 = node1573_r;
      node1576_r = node1464_r & pixel[235];
      node1576_l = node1464_r & ~pixel[235];
      node1577_r = node1576_l & pixel[543];
      node1577_l = node1576_l & ~pixel[543];
      node1578_r = node1577_l & pixel[485];
      node1578_l = node1577_l & ~pixel[485];
      node1579_r = node1578_l & pixel[192];
      node1579_l = node1578_l & ~pixel[192];
      node1580_r = node1579_l & pixel[317];
      node1580_l = node1579_l & ~pixel[317];
      node1581_r = node1580_l & pixel[584];
      node1581_l = node1580_l & ~pixel[584];
      node1582 = node1581_l;
      node1583 = node1581_r;
      node1584_r = node1580_r & pixel[232];
      node1584_l = node1580_r & ~pixel[232];
      node1585 = node1584_l;
      node1586 = node1584_r;
      node1587_r = node1579_r & pixel[321];
      node1587_l = node1579_r & ~pixel[321];
      node1588 = node1587_l;
      node1589_r = node1587_r & pixel[461];
      node1589_l = node1587_r & ~pixel[461];
      node1590 = node1589_l;
      node1591 = node1589_r;
      node1592_r = node1578_r & pixel[289];
      node1592_l = node1578_r & ~pixel[289];
      node1593_r = node1592_l & pixel[551];
      node1593_l = node1592_l & ~pixel[551];
      node1594_r = node1593_l & pixel[292];
      node1594_l = node1593_l & ~pixel[292];
      node1595 = node1594_l;
      node1596 = node1594_r;
      node1597_r = node1593_r & pixel[321];
      node1597_l = node1593_r & ~pixel[321];
      node1598 = node1597_l;
      node1599 = node1597_r;
      node1600_r = node1592_r & pixel[431];
      node1600_l = node1592_r & ~pixel[431];
      node1601_r = node1600_l & pixel[685];
      node1601_l = node1600_l & ~pixel[685];
      node1602 = node1601_l;
      node1603 = node1601_r;
      node1604_r = node1600_r & pixel[159];
      node1604_l = node1600_r & ~pixel[159];
      node1605 = node1604_l;
      node1606 = node1604_r;
      node1607_r = node1577_r & pixel[484];
      node1607_l = node1577_r & ~pixel[484];
      node1608_r = node1607_l & pixel[538];
      node1608_l = node1607_l & ~pixel[538];
      node1609_r = node1608_l & pixel[655];
      node1609_l = node1608_l & ~pixel[655];
      node1610_r = node1609_l & pixel[540];
      node1610_l = node1609_l & ~pixel[540];
      node1611 = node1610_l;
      node1612 = node1610_r;
      node1613_r = node1609_r & pixel[433];
      node1613_l = node1609_r & ~pixel[433];
      node1614 = node1613_l;
      node1615 = node1613_r;
      node1616_r = node1608_r & pixel[599];
      node1616_l = node1608_r & ~pixel[599];
      node1617 = node1616_l;
      node1618_r = node1616_r & pixel[210];
      node1618_l = node1616_r & ~pixel[210];
      node1619 = node1618_l;
      node1620 = node1618_r;
      node1621_r = node1607_r & pixel[479];
      node1621_l = node1607_r & ~pixel[479];
      node1622_r = node1621_l & pixel[554];
      node1622_l = node1621_l & ~pixel[554];
      node1623_r = node1622_l & pixel[411];
      node1623_l = node1622_l & ~pixel[411];
      node1624 = node1623_l;
      node1625 = node1623_r;
      node1626_r = node1622_r & pixel[567];
      node1626_l = node1622_r & ~pixel[567];
      node1627 = node1626_l;
      node1628 = node1626_r;
      node1629 = node1621_r;
      node1630_r = node1576_r & pixel[319];
      node1630_l = node1576_r & ~pixel[319];
      node1631_r = node1630_l & pixel[485];
      node1631_l = node1630_l & ~pixel[485];
      node1632_r = node1631_l & pixel[398];
      node1632_l = node1631_l & ~pixel[398];
      node1633_r = node1632_l & pixel[377];
      node1633_l = node1632_l & ~pixel[377];
      node1634_r = node1633_l & pixel[428];
      node1634_l = node1633_l & ~pixel[428];
      node1635 = node1634_l;
      node1636 = node1634_r;
      node1637_r = node1633_r & pixel[192];
      node1637_l = node1633_r & ~pixel[192];
      node1638 = node1637_l;
      node1639 = node1637_r;
      node1640_r = node1632_r & pixel[634];
      node1640_l = node1632_r & ~pixel[634];
      node1641_r = node1640_l & pixel[429];
      node1641_l = node1640_l & ~pixel[429];
      node1642 = node1641_l;
      node1643 = node1641_r;
      node1644_r = node1640_r & pixel[324];
      node1644_l = node1640_r & ~pixel[324];
      node1645 = node1644_l;
      node1646 = node1644_r;
      node1647_r = node1631_r & pixel[546];
      node1647_l = node1631_r & ~pixel[546];
      node1648_r = node1647_l & pixel[343];
      node1648_l = node1647_l & ~pixel[343];
      node1649_r = node1648_l & pixel[316];
      node1649_l = node1648_l & ~pixel[316];
      node1650 = node1649_l;
      node1651 = node1649_r;
      node1652_r = node1648_r & pixel[101];
      node1652_l = node1648_r & ~pixel[101];
      node1653 = node1652_l;
      node1654 = node1652_r;
      node1655_r = node1647_r & pixel[683];
      node1655_l = node1647_r & ~pixel[683];
      node1656_r = node1655_l & pixel[384];
      node1656_l = node1655_l & ~pixel[384];
      node1657 = node1656_l;
      node1658 = node1656_r;
      node1659_r = node1655_r & pixel[428];
      node1659_l = node1655_r & ~pixel[428];
      node1660 = node1659_l;
      node1661 = node1659_r;
      node1662_r = node1630_r & pixel[490];
      node1662_l = node1630_r & ~pixel[490];
      node1663_r = node1662_l & pixel[405];
      node1663_l = node1662_l & ~pixel[405];
      node1664_r = node1663_l & pixel[272];
      node1664_l = node1663_l & ~pixel[272];
      node1665_r = node1664_l & pixel[189];
      node1665_l = node1664_l & ~pixel[189];
      node1666 = node1665_l;
      node1667 = node1665_r;
      node1668_r = node1664_r & pixel[263];
      node1668_l = node1664_r & ~pixel[263];
      node1669 = node1668_l;
      node1670 = node1668_r;
      node1671_r = node1663_r & pixel[400];
      node1671_l = node1663_r & ~pixel[400];
      node1672_r = node1671_l & pixel[290];
      node1672_l = node1671_l & ~pixel[290];
      node1673 = node1672_l;
      node1674 = node1672_r;
      node1675_r = node1671_r & pixel[213];
      node1675_l = node1671_r & ~pixel[213];
      node1676 = node1675_l;
      node1677 = node1675_r;
      node1678_r = node1662_r & pixel[487];
      node1678_l = node1662_r & ~pixel[487];
      node1679_r = node1678_l & pixel[470];
      node1679_l = node1678_l & ~pixel[470];
      node1680_r = node1679_l & pixel[437];
      node1680_l = node1679_l & ~pixel[437];
      node1681 = node1680_l;
      node1682 = node1680_r;
      node1683_r = node1679_r & pixel[123];
      node1683_l = node1679_r & ~pixel[123];
      node1684 = node1683_l;
      node1685 = node1683_r;
      node1686_r = node1678_r & pixel[427];
      node1686_l = node1678_r & ~pixel[427];
      node1687_r = node1686_l & pixel[471];
      node1687_l = node1686_l & ~pixel[471];
      node1688 = node1687_l;
      node1689 = node1687_r;
      node1690_r = node1686_r & pixel[242];
      node1690_l = node1686_r & ~pixel[242];
      node1691 = node1690_l;
      node1692 = node1690_r;
      result0 = node29 | node52 | node80 | node84 | node92 | node107 | node193 | node338 | node343 | node349 | node350 | node361 | node378 | node398 | node401 | node408 | node409 | node488 | node493 | node502 | node504 | node505 | node510 | node513 | node537 | node547 | node557 | node560 | node571 | node572 | node596 | node608 | node617 | node619 | node620 | node623 | node626 | node808 | node820 | node840 | node843 | node845 | node868 | node875 | node877 | node883 | node885 | node889 | node890 | node893 | node905 | node914 | node921 | node955 | node958 | node972 | node981 | node994 | node998 | node1024 | node1027 | node1038 | node1041 | node1045 | node1047 | node1048 | node1052 | node1053 | node1055 | node1056 | node1060 | node1063 | node1087 | node1103 | node1112 | node1127 | node1134 | node1136 | node1137 | node1151 | node1165 | node1166 | node1181 | node1194 | node1207 | node1217 | node1218 | node1221 | node1224 | node1225 | node1236 | node1245 | node1248 | node1249 | node1258 | node1293 | node1296 | node1335 | node1336 | node1344 | node1364 | node1367 | node1402 | node1418 | node1422 | node1445 | node1480 | node1491 | node1502 | node1505 | node1516;
      result1 = node13 | node135 | node138 | node426 | node451 | node524 | node540 | node677 | node773 | node871 | node1270 | node1271 | node1286 | node1347 | node1526 | node1550 | node1567;
      result2 = node17 | node56 | node60 | node63 | node67 | node73 | node76 | node94 | node100 | node113 | node131 | node141 | node154 | node162 | node163 | node177 | node178 | node180 | node210 | node215 | node223 | node226 | node227 | node286 | node321 | node422 | node528 | node554 | node563 | node639 | node642 | node692 | node703 | node748 | node766 | node781 | node809 | node814 | node822 | node826 | node834 | node856 | node867 | node882 | node886 | node898 | node901 | node902 | node907 | node911 | node922 | node928 | node929 | node932 | node935 | node938 | node939 | node948 | node951 | node966 | node970 | node973 | node1012 | node1016 | node1021 | node1040 | node1072 | node1075 | node1078 | node1086 | node1093 | node1094 | node1109 | node1120 | node1124 | node1128 | node1148 | node1190 | node1193 | node1196 | node1209 | node1241 | node1253 | node1280 | node1308 | node1309 | node1348 | node1350 | node1356 | node1360 | node1385 | node1388 | node1389 | node1395 | node1400 | node1409 | node1415 | node1421 | node1448 | node1449 | node1459 | node1462 | node1463 | node1476 | node1483 | node1488 | node1509 | node1513 | node1522 | node1530 | node1544 | node1553 | node1583 | node1598 | node1612 | node1617 | node1624 | node1627 | node1628 | node1636 | node1643 | node1657 | node1658 | node1685 | node1689 | node1692;
      result3 = node10 | node14 | node21 | node26 | node42 | node51 | node57 | node74 | node77 | node88 | node89 | node95 | node123 | node134 | node147 | node153 | node169 | node173 | node186 | node200 | node229 | node232 | node307 | node312 | node319 | node322 | node327 | node352 | node353 | node364 | node396 | node406 | node429 | node460 | node467 | node544 | node695 | node699 | node712 | node731 | node758 | node765 | node833 | node870 | node899 | node912 | node919 | node984 | node988 | node989 | node993 | node1105 | node1125 | node1278 | node1302 | node1304 | node1305 | node1311 | node1316 | node1332 | node1340 | node1343 | node1351 | node1386 | node1393 | node1401 | node1406 | node1428 | node1435 | node1436 | node1439 | node1443 | node1444 | node1452 | node1457 | node1461 | node1472 | node1475 | node1484 | node1487 | node1498 | node1501 | node1523 | node1529 | node1532 | node1540 | node1543 | node1582 | node1585 | node1591 | node1599 | node1602 | node1611 | node1614 | node1619 | node1620 | node1625 | node1629 | node1638 | node1646 | node1650 | node1661 | node1669 | node1673 | node1682;
      result4 = node25 | node36 | node41 | node49 | node83 | node103 | node132 | node139 | node149 | node165 | node195 | node199 | node203 | node207 | node208 | node217 | node243 | node262 | node270 | node273 | node280 | node281 | node288 | node289 | node296 | node297 | node314 | node337 | node367 | node371 | node376 | node383 | node385 | node386 | node391 | node393 | node405 | node444 | node452 | node475 | node478 | node481 | node482 | node490 | node517 | node525 | node556 | node561 | node568 | node650 | node653 | node658 | node667 | node670 | node671 | node685 | node728 | node734 | node797 | node805 | node829 | node832 | node851 | node1152 | node1158 | node1244 | node1273 | node1274 | node1292 | node1357 | node1378 | node1408 | node1559 | node1572;
      result5 = node28 | node35 | node81 | node121 | node142 | node202 | node231 | node246 | node255 | node265 | node266 | node285 | node300 | node303 | node306 | node330 | node331 | node335 | node342 | node345 | node363 | node402 | node430 | node447 | node459 | node487 | node545 | node564 | node579 | node585 | node588 | node603 | node610 | node611 | node616 | node624 | node627 | node660 | node664 | node684 | node687 | node709 | node716 | node717 | node719 | node740 | node751 | node755 | node756 | node780 | node783 | node874 | node915 | node918 | node931 | node947 | node962 | node969 | node980 | node983 | node987 | node995 | node1005 | node1008 | node1020 | node1031 | node1044 | node1062 | node1068 | node1076 | node1102 | node1106 | node1133 | node1141 | node1143 | node1144 | node1167 | node1168 | node1172 | node1176 | node1201 | node1210 | node1227 | node1237 | node1281 | node1289 | node1317 | node1319 | node1320 | node1331 | node1334 | node1392 | node1431 | node1438 | node1471 | node1481 | node1490 | node1496 | node1497 | node1504 | node1515 | node1564 | node1571 | node1586 | node1588 | node1590 | node1603 | node1639 | node1645 | node1666 | node1667 | node1670 | node1677;
      result6 = node11 | node32 | node33 | node45 | node48 | node64 | node66 | node101 | node104 | node108 | node109 | node114 | node116 | node124 | node157 | node166 | node181 | node192 | node211 | node214 | node218 | node237 | node244 | node282 | node290 | node328 | node334 | node368 | node382 | node392 | node397 | node410 | node435 | node438 | node439 | node454 | node461 | node491 | node495 | node496 | node506 | node516 | node527 | node548 | node553 | node569 | node578 | node634 | node635 | node654 | node702 | node747 | node774 | node776 | node777 | node785 | node790 | node791 | node794 | node801 | node806 | node828 | node838 | node841 | node846 | node854 | node892 | node950 | node963 | node965 | node1023 | node1028 | node1030 | node1037 | node1071 | node1083 | node1084 | node1091 | node1113 | node1121 | node1173 | node1175 | node1179 | node1186 | node1187 | node1189 | node1197 | node1228 | node1229 | node1230 | node1235 | node1242 | node1260 | node1295 | node1325 | node1363 | node1366 | node1405 | node1414 | node1417 | node1525 | node1533 | node1556 | node1642 | node1654 | node1676 | node1684 | node1691;
      result7 = node18 | node44 | node146 | node185 | node256 | node258 | node263 | node271 | node275 | node360 | node379 | node419 | node420 | node423 | node434 | node464 | node474 | node501 | node509 | node531 | node541 | node592 | node600 | node607 | node680 | node700 | node735 | node941 | node1117 | node1155 | node1250 | node1288 | node1370 | node1374 | node1377;
      result8 = node20 | node90 | node117 | node150 | node156 | node240 | node247 | node259 | node274 | node304 | node315 | node318 | node346 | node370 | node427 | node455 | node532 | node538 | node576 | node632 | node641 | node666 | node672 | node710 | node713 | node720 | node725 | node741 | node743 | node744 | node762 | node763 | node784 | node793 | node798 | node812 | node813 | node821 | node825 | node849 | node857 | node878 | node906 | node936 | node954 | node957 | node999 | node1006 | node1009 | node1013 | node1015 | node1059 | node1069 | node1079 | node1090 | node1110 | node1118 | node1140 | node1149 | node1159 | node1180 | node1202 | node1203 | node1206 | node1254 | node1261 | node1277 | node1285 | node1301 | node1312 | node1323 | node1324 | node1341 | node1359 | node1371 | node1375 | node1396 | node1419 | node1429 | node1432 | node1451 | node1456 | node1474 | node1511 | node1537 | node1538 | node1541 | node1549 | node1552 | node1557 | node1560 | node1565 | node1568 | node1574 | node1575 | node1595 | node1596 | node1605 | node1606 | node1615 | node1635 | node1651 | node1653 | node1660 | node1674 | node1681 | node1688;
      result9 = node59 | node120 | node170 | node172 | node183 | node196 | node224 | node236 | node239 | node299 | node311 | node375 | node437 | node445 | node448 | node465 | node468 | node477 | node483 | node514 | node533 | node575 | node586 | node589 | node593 | node595 | node601 | node604 | node631 | node638 | node651 | node657 | node661 | node678 | node681 | node688 | node693 | node696 | node724 | node727 | node732 | node750 | node759 | node800 | node852 | node942 | node1000 | node1156 | node1220 | node1257 | node1510;

      tree_0 = {result9, result8, result7, result6, result5, result4, result3, result2, result1, result0};
    end
  endfunction

  function [9:0] tree_1;
    input [783:0] pixel;

    reg node0_r;
    reg node0_l;
    reg node1_r;
    reg node1_l;
    reg node2_r;
    reg node2_l;
    reg node3_r;
    reg node3_l;
    reg node4_r;
    reg node4_l;
    reg node5_r;
    reg node5_l;
    reg node6_r;
    reg node6_l;
    reg node7_r;
    reg node7_l;
    reg node8_r;
    reg node8_l;
    reg node9_r;
    reg node9_l;
    reg node10;
    reg node11;
    reg node12_r;
    reg node12_l;
    reg node13;
    reg node14;
    reg node15_r;
    reg node15_l;
    reg node16_r;
    reg node16_l;
    reg node17;
    reg node18;
    reg node19_r;
    reg node19_l;
    reg node20;
    reg node21;
    reg node22_r;
    reg node22_l;
    reg node23_r;
    reg node23_l;
    reg node24;
    reg node25;
    reg node26;
    reg node27_r;
    reg node27_l;
    reg node28_r;
    reg node28_l;
    reg node29_r;
    reg node29_l;
    reg node30_r;
    reg node30_l;
    reg node31;
    reg node32;
    reg node33_r;
    reg node33_l;
    reg node34;
    reg node35;
    reg node36_r;
    reg node36_l;
    reg node37_r;
    reg node37_l;
    reg node38;
    reg node39;
    reg node40_r;
    reg node40_l;
    reg node41;
    reg node42;
    reg node43_r;
    reg node43_l;
    reg node44_r;
    reg node44_l;
    reg node45_r;
    reg node45_l;
    reg node46;
    reg node47;
    reg node48_r;
    reg node48_l;
    reg node49;
    reg node50;
    reg node51_r;
    reg node51_l;
    reg node52_r;
    reg node52_l;
    reg node53;
    reg node54;
    reg node55_r;
    reg node55_l;
    reg node56;
    reg node57;
    reg node58_r;
    reg node58_l;
    reg node59_r;
    reg node59_l;
    reg node60_r;
    reg node60_l;
    reg node61_r;
    reg node61_l;
    reg node62_r;
    reg node62_l;
    reg node63;
    reg node64;
    reg node65_r;
    reg node65_l;
    reg node66;
    reg node67;
    reg node68_r;
    reg node68_l;
    reg node69;
    reg node70;
    reg node71_r;
    reg node71_l;
    reg node72_r;
    reg node72_l;
    reg node73;
    reg node74_r;
    reg node74_l;
    reg node75;
    reg node76;
    reg node77_r;
    reg node77_l;
    reg node78;
    reg node79;
    reg node80_r;
    reg node80_l;
    reg node81_r;
    reg node81_l;
    reg node82_r;
    reg node82_l;
    reg node83_r;
    reg node83_l;
    reg node84;
    reg node85;
    reg node86;
    reg node87_r;
    reg node87_l;
    reg node88_r;
    reg node88_l;
    reg node89;
    reg node90;
    reg node91;
    reg node92_r;
    reg node92_l;
    reg node93;
    reg node94;
    reg node95_r;
    reg node95_l;
    reg node96_r;
    reg node96_l;
    reg node97_r;
    reg node97_l;
    reg node98_r;
    reg node98_l;
    reg node99_r;
    reg node99_l;
    reg node100_r;
    reg node100_l;
    reg node101;
    reg node102;
    reg node103;
    reg node104_r;
    reg node104_l;
    reg node105_r;
    reg node105_l;
    reg node106;
    reg node107;
    reg node108;
    reg node109_r;
    reg node109_l;
    reg node110_r;
    reg node110_l;
    reg node111_r;
    reg node111_l;
    reg node112;
    reg node113;
    reg node114_r;
    reg node114_l;
    reg node115;
    reg node116;
    reg node117_r;
    reg node117_l;
    reg node118_r;
    reg node118_l;
    reg node119;
    reg node120;
    reg node121;
    reg node122_r;
    reg node122_l;
    reg node123_r;
    reg node123_l;
    reg node124_r;
    reg node124_l;
    reg node125_r;
    reg node125_l;
    reg node126;
    reg node127;
    reg node128_r;
    reg node128_l;
    reg node129;
    reg node130;
    reg node131_r;
    reg node131_l;
    reg node132_r;
    reg node132_l;
    reg node133;
    reg node134;
    reg node135_r;
    reg node135_l;
    reg node136;
    reg node137;
    reg node138_r;
    reg node138_l;
    reg node139_r;
    reg node139_l;
    reg node140_r;
    reg node140_l;
    reg node141;
    reg node142;
    reg node143_r;
    reg node143_l;
    reg node144;
    reg node145;
    reg node146_r;
    reg node146_l;
    reg node147_r;
    reg node147_l;
    reg node148;
    reg node149;
    reg node150_r;
    reg node150_l;
    reg node151;
    reg node152;
    reg node153_r;
    reg node153_l;
    reg node154_r;
    reg node154_l;
    reg node155_r;
    reg node155_l;
    reg node156_r;
    reg node156_l;
    reg node157_r;
    reg node157_l;
    reg node158;
    reg node159;
    reg node160_r;
    reg node160_l;
    reg node161;
    reg node162;
    reg node163_r;
    reg node163_l;
    reg node164_r;
    reg node164_l;
    reg node165;
    reg node166;
    reg node167_r;
    reg node167_l;
    reg node168;
    reg node169;
    reg node170_r;
    reg node170_l;
    reg node171_r;
    reg node171_l;
    reg node172_r;
    reg node172_l;
    reg node173;
    reg node174;
    reg node175;
    reg node176_r;
    reg node176_l;
    reg node177;
    reg node178;
    reg node179_r;
    reg node179_l;
    reg node180_r;
    reg node180_l;
    reg node181_r;
    reg node181_l;
    reg node182_r;
    reg node182_l;
    reg node183;
    reg node184;
    reg node185;
    reg node186_r;
    reg node186_l;
    reg node187;
    reg node188_r;
    reg node188_l;
    reg node189;
    reg node190;
    reg node191_r;
    reg node191_l;
    reg node192_r;
    reg node192_l;
    reg node193_r;
    reg node193_l;
    reg node194;
    reg node195;
    reg node196_r;
    reg node196_l;
    reg node197;
    reg node198;
    reg node199_r;
    reg node199_l;
    reg node200;
    reg node201_r;
    reg node201_l;
    reg node202;
    reg node203;
    reg node204_r;
    reg node204_l;
    reg node205_r;
    reg node205_l;
    reg node206_r;
    reg node206_l;
    reg node207_r;
    reg node207_l;
    reg node208_r;
    reg node208_l;
    reg node209_r;
    reg node209_l;
    reg node210_r;
    reg node210_l;
    reg node211;
    reg node212;
    reg node213_r;
    reg node213_l;
    reg node214;
    reg node215;
    reg node216_r;
    reg node216_l;
    reg node217_r;
    reg node217_l;
    reg node218;
    reg node219;
    reg node220;
    reg node221_r;
    reg node221_l;
    reg node222_r;
    reg node222_l;
    reg node223_r;
    reg node223_l;
    reg node224;
    reg node225;
    reg node226_r;
    reg node226_l;
    reg node227;
    reg node228;
    reg node229_r;
    reg node229_l;
    reg node230_r;
    reg node230_l;
    reg node231;
    reg node232;
    reg node233_r;
    reg node233_l;
    reg node234;
    reg node235;
    reg node236_r;
    reg node236_l;
    reg node237_r;
    reg node237_l;
    reg node238_r;
    reg node238_l;
    reg node239_r;
    reg node239_l;
    reg node240;
    reg node241;
    reg node242_r;
    reg node242_l;
    reg node243;
    reg node244;
    reg node245_r;
    reg node245_l;
    reg node246_r;
    reg node246_l;
    reg node247;
    reg node248;
    reg node249_r;
    reg node249_l;
    reg node250;
    reg node251;
    reg node252_r;
    reg node252_l;
    reg node253_r;
    reg node253_l;
    reg node254_r;
    reg node254_l;
    reg node255;
    reg node256;
    reg node257_r;
    reg node257_l;
    reg node258;
    reg node259;
    reg node260_r;
    reg node260_l;
    reg node261_r;
    reg node261_l;
    reg node262;
    reg node263;
    reg node264;
    reg node265_r;
    reg node265_l;
    reg node266_r;
    reg node266_l;
    reg node267_r;
    reg node267_l;
    reg node268_r;
    reg node268_l;
    reg node269_r;
    reg node269_l;
    reg node270;
    reg node271;
    reg node272_r;
    reg node272_l;
    reg node273;
    reg node274;
    reg node275;
    reg node276_r;
    reg node276_l;
    reg node277_r;
    reg node277_l;
    reg node278_r;
    reg node278_l;
    reg node279;
    reg node280;
    reg node281_r;
    reg node281_l;
    reg node282;
    reg node283;
    reg node284_r;
    reg node284_l;
    reg node285_r;
    reg node285_l;
    reg node286;
    reg node287;
    reg node288_r;
    reg node288_l;
    reg node289;
    reg node290;
    reg node291_r;
    reg node291_l;
    reg node292_r;
    reg node292_l;
    reg node293_r;
    reg node293_l;
    reg node294_r;
    reg node294_l;
    reg node295;
    reg node296;
    reg node297_r;
    reg node297_l;
    reg node298;
    reg node299;
    reg node300_r;
    reg node300_l;
    reg node301_r;
    reg node301_l;
    reg node302;
    reg node303;
    reg node304;
    reg node305_r;
    reg node305_l;
    reg node306_r;
    reg node306_l;
    reg node307_r;
    reg node307_l;
    reg node308;
    reg node309;
    reg node310_r;
    reg node310_l;
    reg node311;
    reg node312;
    reg node313_r;
    reg node313_l;
    reg node314_r;
    reg node314_l;
    reg node315;
    reg node316;
    reg node317_r;
    reg node317_l;
    reg node318;
    reg node319;
    reg node320_r;
    reg node320_l;
    reg node321_r;
    reg node321_l;
    reg node322_r;
    reg node322_l;
    reg node323_r;
    reg node323_l;
    reg node324_r;
    reg node324_l;
    reg node325_r;
    reg node325_l;
    reg node326;
    reg node327;
    reg node328_r;
    reg node328_l;
    reg node329;
    reg node330;
    reg node331_r;
    reg node331_l;
    reg node332_r;
    reg node332_l;
    reg node333;
    reg node334;
    reg node335;
    reg node336_r;
    reg node336_l;
    reg node337_r;
    reg node337_l;
    reg node338_r;
    reg node338_l;
    reg node339;
    reg node340;
    reg node341_r;
    reg node341_l;
    reg node342;
    reg node343;
    reg node344_r;
    reg node344_l;
    reg node345_r;
    reg node345_l;
    reg node346;
    reg node347;
    reg node348_r;
    reg node348_l;
    reg node349;
    reg node350;
    reg node351_r;
    reg node351_l;
    reg node352_r;
    reg node352_l;
    reg node353_r;
    reg node353_l;
    reg node354_r;
    reg node354_l;
    reg node355;
    reg node356;
    reg node357_r;
    reg node357_l;
    reg node358;
    reg node359;
    reg node360_r;
    reg node360_l;
    reg node361_r;
    reg node361_l;
    reg node362;
    reg node363;
    reg node364_r;
    reg node364_l;
    reg node365;
    reg node366;
    reg node367_r;
    reg node367_l;
    reg node368_r;
    reg node368_l;
    reg node369_r;
    reg node369_l;
    reg node370;
    reg node371;
    reg node372_r;
    reg node372_l;
    reg node373;
    reg node374;
    reg node375_r;
    reg node375_l;
    reg node376_r;
    reg node376_l;
    reg node377;
    reg node378;
    reg node379_r;
    reg node379_l;
    reg node380;
    reg node381;
    reg node382_r;
    reg node382_l;
    reg node383_r;
    reg node383_l;
    reg node384_r;
    reg node384_l;
    reg node385_r;
    reg node385_l;
    reg node386_r;
    reg node386_l;
    reg node387;
    reg node388;
    reg node389_r;
    reg node389_l;
    reg node390;
    reg node391;
    reg node392_r;
    reg node392_l;
    reg node393_r;
    reg node393_l;
    reg node394;
    reg node395;
    reg node396_r;
    reg node396_l;
    reg node397;
    reg node398;
    reg node399_r;
    reg node399_l;
    reg node400_r;
    reg node400_l;
    reg node401_r;
    reg node401_l;
    reg node402;
    reg node403;
    reg node404;
    reg node405;
    reg node406_r;
    reg node406_l;
    reg node407_r;
    reg node407_l;
    reg node408_r;
    reg node408_l;
    reg node409_r;
    reg node409_l;
    reg node410;
    reg node411;
    reg node412_r;
    reg node412_l;
    reg node413;
    reg node414;
    reg node415_r;
    reg node415_l;
    reg node416;
    reg node417;
    reg node418_r;
    reg node418_l;
    reg node419_r;
    reg node419_l;
    reg node420_r;
    reg node420_l;
    reg node421;
    reg node422;
    reg node423;
    reg node424_r;
    reg node424_l;
    reg node425;
    reg node426;
    reg node427_r;
    reg node427_l;
    reg node428_r;
    reg node428_l;
    reg node429_r;
    reg node429_l;
    reg node430_r;
    reg node430_l;
    reg node431_r;
    reg node431_l;
    reg node432_r;
    reg node432_l;
    reg node433_r;
    reg node433_l;
    reg node434_r;
    reg node434_l;
    reg node435;
    reg node436;
    reg node437_r;
    reg node437_l;
    reg node438;
    reg node439;
    reg node440_r;
    reg node440_l;
    reg node441_r;
    reg node441_l;
    reg node442;
    reg node443;
    reg node444_r;
    reg node444_l;
    reg node445;
    reg node446;
    reg node447_r;
    reg node447_l;
    reg node448_r;
    reg node448_l;
    reg node449_r;
    reg node449_l;
    reg node450;
    reg node451;
    reg node452_r;
    reg node452_l;
    reg node453;
    reg node454;
    reg node455_r;
    reg node455_l;
    reg node456_r;
    reg node456_l;
    reg node457;
    reg node458;
    reg node459_r;
    reg node459_l;
    reg node460;
    reg node461;
    reg node462_r;
    reg node462_l;
    reg node463_r;
    reg node463_l;
    reg node464_r;
    reg node464_l;
    reg node465_r;
    reg node465_l;
    reg node466;
    reg node467;
    reg node468_r;
    reg node468_l;
    reg node469;
    reg node470;
    reg node471_r;
    reg node471_l;
    reg node472_r;
    reg node472_l;
    reg node473;
    reg node474;
    reg node475_r;
    reg node475_l;
    reg node476;
    reg node477;
    reg node478_r;
    reg node478_l;
    reg node479_r;
    reg node479_l;
    reg node480_r;
    reg node480_l;
    reg node481;
    reg node482;
    reg node483_r;
    reg node483_l;
    reg node484;
    reg node485;
    reg node486_r;
    reg node486_l;
    reg node487_r;
    reg node487_l;
    reg node488;
    reg node489;
    reg node490_r;
    reg node490_l;
    reg node491;
    reg node492;
    reg node493_r;
    reg node493_l;
    reg node494_r;
    reg node494_l;
    reg node495_r;
    reg node495_l;
    reg node496_r;
    reg node496_l;
    reg node497_r;
    reg node497_l;
    reg node498;
    reg node499;
    reg node500_r;
    reg node500_l;
    reg node501;
    reg node502;
    reg node503_r;
    reg node503_l;
    reg node504_r;
    reg node504_l;
    reg node505;
    reg node506;
    reg node507_r;
    reg node507_l;
    reg node508;
    reg node509;
    reg node510_r;
    reg node510_l;
    reg node511_r;
    reg node511_l;
    reg node512_r;
    reg node512_l;
    reg node513;
    reg node514;
    reg node515_r;
    reg node515_l;
    reg node516;
    reg node517;
    reg node518_r;
    reg node518_l;
    reg node519_r;
    reg node519_l;
    reg node520;
    reg node521;
    reg node522_r;
    reg node522_l;
    reg node523;
    reg node524;
    reg node525_r;
    reg node525_l;
    reg node526_r;
    reg node526_l;
    reg node527_r;
    reg node527_l;
    reg node528_r;
    reg node528_l;
    reg node529;
    reg node530;
    reg node531;
    reg node532_r;
    reg node532_l;
    reg node533_r;
    reg node533_l;
    reg node534;
    reg node535;
    reg node536_r;
    reg node536_l;
    reg node537;
    reg node538;
    reg node539_r;
    reg node539_l;
    reg node540_r;
    reg node540_l;
    reg node541_r;
    reg node541_l;
    reg node542;
    reg node543;
    reg node544_r;
    reg node544_l;
    reg node545;
    reg node546;
    reg node547_r;
    reg node547_l;
    reg node548_r;
    reg node548_l;
    reg node549;
    reg node550;
    reg node551_r;
    reg node551_l;
    reg node552;
    reg node553;
    reg node554_r;
    reg node554_l;
    reg node555_r;
    reg node555_l;
    reg node556_r;
    reg node556_l;
    reg node557_r;
    reg node557_l;
    reg node558_r;
    reg node558_l;
    reg node559_r;
    reg node559_l;
    reg node560;
    reg node561;
    reg node562_r;
    reg node562_l;
    reg node563;
    reg node564;
    reg node565_r;
    reg node565_l;
    reg node566_r;
    reg node566_l;
    reg node567;
    reg node568;
    reg node569_r;
    reg node569_l;
    reg node570;
    reg node571;
    reg node572_r;
    reg node572_l;
    reg node573_r;
    reg node573_l;
    reg node574_r;
    reg node574_l;
    reg node575;
    reg node576;
    reg node577_r;
    reg node577_l;
    reg node578;
    reg node579;
    reg node580_r;
    reg node580_l;
    reg node581;
    reg node582_r;
    reg node582_l;
    reg node583;
    reg node584;
    reg node585_r;
    reg node585_l;
    reg node586_r;
    reg node586_l;
    reg node587_r;
    reg node587_l;
    reg node588_r;
    reg node588_l;
    reg node589;
    reg node590;
    reg node591;
    reg node592;
    reg node593_r;
    reg node593_l;
    reg node594;
    reg node595_r;
    reg node595_l;
    reg node596;
    reg node597;
    reg node598_r;
    reg node598_l;
    reg node599_r;
    reg node599_l;
    reg node600_r;
    reg node600_l;
    reg node601_r;
    reg node601_l;
    reg node602_r;
    reg node602_l;
    reg node603;
    reg node604;
    reg node605_r;
    reg node605_l;
    reg node606;
    reg node607;
    reg node608_r;
    reg node608_l;
    reg node609_r;
    reg node609_l;
    reg node610;
    reg node611;
    reg node612_r;
    reg node612_l;
    reg node613;
    reg node614;
    reg node615_r;
    reg node615_l;
    reg node616_r;
    reg node616_l;
    reg node617_r;
    reg node617_l;
    reg node618;
    reg node619;
    reg node620_r;
    reg node620_l;
    reg node621;
    reg node622;
    reg node623_r;
    reg node623_l;
    reg node624_r;
    reg node624_l;
    reg node625;
    reg node626;
    reg node627_r;
    reg node627_l;
    reg node628;
    reg node629;
    reg node630_r;
    reg node630_l;
    reg node631_r;
    reg node631_l;
    reg node632_r;
    reg node632_l;
    reg node633_r;
    reg node633_l;
    reg node634;
    reg node635;
    reg node636_r;
    reg node636_l;
    reg node637;
    reg node638;
    reg node639_r;
    reg node639_l;
    reg node640_r;
    reg node640_l;
    reg node641;
    reg node642;
    reg node643_r;
    reg node643_l;
    reg node644;
    reg node645;
    reg node646_r;
    reg node646_l;
    reg node647_r;
    reg node647_l;
    reg node648_r;
    reg node648_l;
    reg node649;
    reg node650;
    reg node651_r;
    reg node651_l;
    reg node652;
    reg node653;
    reg node654_r;
    reg node654_l;
    reg node655_r;
    reg node655_l;
    reg node656;
    reg node657;
    reg node658_r;
    reg node658_l;
    reg node659;
    reg node660;
    reg node661_r;
    reg node661_l;
    reg node662_r;
    reg node662_l;
    reg node663_r;
    reg node663_l;
    reg node664_r;
    reg node664_l;
    reg node665_r;
    reg node665_l;
    reg node666_r;
    reg node666_l;
    reg node667_r;
    reg node667_l;
    reg node668;
    reg node669;
    reg node670_r;
    reg node670_l;
    reg node671;
    reg node672;
    reg node673_r;
    reg node673_l;
    reg node674_r;
    reg node674_l;
    reg node675;
    reg node676;
    reg node677_r;
    reg node677_l;
    reg node678;
    reg node679;
    reg node680_r;
    reg node680_l;
    reg node681_r;
    reg node681_l;
    reg node682_r;
    reg node682_l;
    reg node683;
    reg node684;
    reg node685_r;
    reg node685_l;
    reg node686;
    reg node687;
    reg node688_r;
    reg node688_l;
    reg node689_r;
    reg node689_l;
    reg node690;
    reg node691;
    reg node692_r;
    reg node692_l;
    reg node693;
    reg node694;
    reg node695_r;
    reg node695_l;
    reg node696_r;
    reg node696_l;
    reg node697_r;
    reg node697_l;
    reg node698_r;
    reg node698_l;
    reg node699;
    reg node700;
    reg node701_r;
    reg node701_l;
    reg node702;
    reg node703;
    reg node704_r;
    reg node704_l;
    reg node705_r;
    reg node705_l;
    reg node706;
    reg node707;
    reg node708_r;
    reg node708_l;
    reg node709;
    reg node710;
    reg node711_r;
    reg node711_l;
    reg node712_r;
    reg node712_l;
    reg node713_r;
    reg node713_l;
    reg node714;
    reg node715;
    reg node716_r;
    reg node716_l;
    reg node717;
    reg node718;
    reg node719_r;
    reg node719_l;
    reg node720_r;
    reg node720_l;
    reg node721;
    reg node722;
    reg node723_r;
    reg node723_l;
    reg node724;
    reg node725;
    reg node726_r;
    reg node726_l;
    reg node727_r;
    reg node727_l;
    reg node728_r;
    reg node728_l;
    reg node729_r;
    reg node729_l;
    reg node730;
    reg node731_r;
    reg node731_l;
    reg node732;
    reg node733;
    reg node734_r;
    reg node734_l;
    reg node735_r;
    reg node735_l;
    reg node736;
    reg node737;
    reg node738_r;
    reg node738_l;
    reg node739;
    reg node740;
    reg node741_r;
    reg node741_l;
    reg node742_r;
    reg node742_l;
    reg node743_r;
    reg node743_l;
    reg node744;
    reg node745;
    reg node746_r;
    reg node746_l;
    reg node747;
    reg node748;
    reg node749_r;
    reg node749_l;
    reg node750_r;
    reg node750_l;
    reg node751;
    reg node752;
    reg node753_r;
    reg node753_l;
    reg node754;
    reg node755;
    reg node756_r;
    reg node756_l;
    reg node757_r;
    reg node757_l;
    reg node758_r;
    reg node758_l;
    reg node759_r;
    reg node759_l;
    reg node760;
    reg node761;
    reg node762_r;
    reg node762_l;
    reg node763;
    reg node764;
    reg node765_r;
    reg node765_l;
    reg node766_r;
    reg node766_l;
    reg node767;
    reg node768;
    reg node769_r;
    reg node769_l;
    reg node770;
    reg node771;
    reg node772_r;
    reg node772_l;
    reg node773_r;
    reg node773_l;
    reg node774_r;
    reg node774_l;
    reg node775;
    reg node776;
    reg node777;
    reg node778;
    reg node779_r;
    reg node779_l;
    reg node780_r;
    reg node780_l;
    reg node781_r;
    reg node781_l;
    reg node782_r;
    reg node782_l;
    reg node783_r;
    reg node783_l;
    reg node784;
    reg node785_r;
    reg node785_l;
    reg node786;
    reg node787;
    reg node788_r;
    reg node788_l;
    reg node789_r;
    reg node789_l;
    reg node790;
    reg node791;
    reg node792_r;
    reg node792_l;
    reg node793;
    reg node794;
    reg node795_r;
    reg node795_l;
    reg node796;
    reg node797_r;
    reg node797_l;
    reg node798_r;
    reg node798_l;
    reg node799;
    reg node800;
    reg node801_r;
    reg node801_l;
    reg node802;
    reg node803;
    reg node804_r;
    reg node804_l;
    reg node805_r;
    reg node805_l;
    reg node806_r;
    reg node806_l;
    reg node807_r;
    reg node807_l;
    reg node808;
    reg node809;
    reg node810;
    reg node811_r;
    reg node811_l;
    reg node812_r;
    reg node812_l;
    reg node813;
    reg node814;
    reg node815_r;
    reg node815_l;
    reg node816;
    reg node817;
    reg node818_r;
    reg node818_l;
    reg node819_r;
    reg node819_l;
    reg node820_r;
    reg node820_l;
    reg node821;
    reg node822;
    reg node823_r;
    reg node823_l;
    reg node824;
    reg node825;
    reg node826_r;
    reg node826_l;
    reg node827_r;
    reg node827_l;
    reg node828;
    reg node829;
    reg node830_r;
    reg node830_l;
    reg node831;
    reg node832;
    reg node833_r;
    reg node833_l;
    reg node834_r;
    reg node834_l;
    reg node835_r;
    reg node835_l;
    reg node836_r;
    reg node836_l;
    reg node837_r;
    reg node837_l;
    reg node838;
    reg node839;
    reg node840_r;
    reg node840_l;
    reg node841;
    reg node842;
    reg node843_r;
    reg node843_l;
    reg node844;
    reg node845_r;
    reg node845_l;
    reg node846;
    reg node847;
    reg node848_r;
    reg node848_l;
    reg node849_r;
    reg node849_l;
    reg node850_r;
    reg node850_l;
    reg node851;
    reg node852;
    reg node853_r;
    reg node853_l;
    reg node854;
    reg node855;
    reg node856_r;
    reg node856_l;
    reg node857_r;
    reg node857_l;
    reg node858;
    reg node859;
    reg node860_r;
    reg node860_l;
    reg node861;
    reg node862;
    reg node863_r;
    reg node863_l;
    reg node864_r;
    reg node864_l;
    reg node865;
    reg node866;
    reg node867_r;
    reg node867_l;
    reg node868_r;
    reg node868_l;
    reg node869;
    reg node870_r;
    reg node870_l;
    reg node871;
    reg node872;
    reg node873_r;
    reg node873_l;
    reg node874_r;
    reg node874_l;
    reg node875;
    reg node876;
    reg node877_r;
    reg node877_l;
    reg node878;
    reg node879;
    reg node880_r;
    reg node880_l;
    reg node881_r;
    reg node881_l;
    reg node882_r;
    reg node882_l;
    reg node883_r;
    reg node883_l;
    reg node884_r;
    reg node884_l;
    reg node885_r;
    reg node885_l;
    reg node886_r;
    reg node886_l;
    reg node887_r;
    reg node887_l;
    reg node888_r;
    reg node888_l;
    reg node889;
    reg node890;
    reg node891_r;
    reg node891_l;
    reg node892;
    reg node893;
    reg node894_r;
    reg node894_l;
    reg node895_r;
    reg node895_l;
    reg node896;
    reg node897;
    reg node898_r;
    reg node898_l;
    reg node899;
    reg node900;
    reg node901_r;
    reg node901_l;
    reg node902_r;
    reg node902_l;
    reg node903_r;
    reg node903_l;
    reg node904;
    reg node905;
    reg node906_r;
    reg node906_l;
    reg node907;
    reg node908;
    reg node909_r;
    reg node909_l;
    reg node910_r;
    reg node910_l;
    reg node911;
    reg node912;
    reg node913_r;
    reg node913_l;
    reg node914;
    reg node915;
    reg node916_r;
    reg node916_l;
    reg node917_r;
    reg node917_l;
    reg node918_r;
    reg node918_l;
    reg node919_r;
    reg node919_l;
    reg node920;
    reg node921;
    reg node922_r;
    reg node922_l;
    reg node923;
    reg node924;
    reg node925_r;
    reg node925_l;
    reg node926_r;
    reg node926_l;
    reg node927;
    reg node928;
    reg node929_r;
    reg node929_l;
    reg node930;
    reg node931;
    reg node932_r;
    reg node932_l;
    reg node933_r;
    reg node933_l;
    reg node934_r;
    reg node934_l;
    reg node935;
    reg node936;
    reg node937_r;
    reg node937_l;
    reg node938;
    reg node939;
    reg node940_r;
    reg node940_l;
    reg node941_r;
    reg node941_l;
    reg node942;
    reg node943;
    reg node944_r;
    reg node944_l;
    reg node945;
    reg node946;
    reg node947_r;
    reg node947_l;
    reg node948_r;
    reg node948_l;
    reg node949_r;
    reg node949_l;
    reg node950_r;
    reg node950_l;
    reg node951_r;
    reg node951_l;
    reg node952;
    reg node953;
    reg node954_r;
    reg node954_l;
    reg node955;
    reg node956;
    reg node957_r;
    reg node957_l;
    reg node958_r;
    reg node958_l;
    reg node959;
    reg node960;
    reg node961_r;
    reg node961_l;
    reg node962;
    reg node963;
    reg node964_r;
    reg node964_l;
    reg node965_r;
    reg node965_l;
    reg node966_r;
    reg node966_l;
    reg node967;
    reg node968;
    reg node969_r;
    reg node969_l;
    reg node970;
    reg node971;
    reg node972;
    reg node973_r;
    reg node973_l;
    reg node974_r;
    reg node974_l;
    reg node975_r;
    reg node975_l;
    reg node976_r;
    reg node976_l;
    reg node977;
    reg node978;
    reg node979_r;
    reg node979_l;
    reg node980;
    reg node981;
    reg node982_r;
    reg node982_l;
    reg node983_r;
    reg node983_l;
    reg node984;
    reg node985;
    reg node986_r;
    reg node986_l;
    reg node987;
    reg node988;
    reg node989_r;
    reg node989_l;
    reg node990_r;
    reg node990_l;
    reg node991_r;
    reg node991_l;
    reg node992;
    reg node993;
    reg node994;
    reg node995;
    reg node996_r;
    reg node996_l;
    reg node997_r;
    reg node997_l;
    reg node998_r;
    reg node998_l;
    reg node999_r;
    reg node999_l;
    reg node1000_r;
    reg node1000_l;
    reg node1001_r;
    reg node1001_l;
    reg node1002;
    reg node1003;
    reg node1004_r;
    reg node1004_l;
    reg node1005;
    reg node1006;
    reg node1007_r;
    reg node1007_l;
    reg node1008_r;
    reg node1008_l;
    reg node1009;
    reg node1010;
    reg node1011_r;
    reg node1011_l;
    reg node1012;
    reg node1013;
    reg node1014_r;
    reg node1014_l;
    reg node1015_r;
    reg node1015_l;
    reg node1016_r;
    reg node1016_l;
    reg node1017;
    reg node1018;
    reg node1019_r;
    reg node1019_l;
    reg node1020;
    reg node1021;
    reg node1022_r;
    reg node1022_l;
    reg node1023_r;
    reg node1023_l;
    reg node1024;
    reg node1025;
    reg node1026_r;
    reg node1026_l;
    reg node1027;
    reg node1028;
    reg node1029_r;
    reg node1029_l;
    reg node1030_r;
    reg node1030_l;
    reg node1031_r;
    reg node1031_l;
    reg node1032_r;
    reg node1032_l;
    reg node1033;
    reg node1034;
    reg node1035_r;
    reg node1035_l;
    reg node1036;
    reg node1037;
    reg node1038_r;
    reg node1038_l;
    reg node1039_r;
    reg node1039_l;
    reg node1040;
    reg node1041;
    reg node1042_r;
    reg node1042_l;
    reg node1043;
    reg node1044;
    reg node1045_r;
    reg node1045_l;
    reg node1046_r;
    reg node1046_l;
    reg node1047_r;
    reg node1047_l;
    reg node1048;
    reg node1049;
    reg node1050_r;
    reg node1050_l;
    reg node1051;
    reg node1052;
    reg node1053_r;
    reg node1053_l;
    reg node1054_r;
    reg node1054_l;
    reg node1055;
    reg node1056;
    reg node1057_r;
    reg node1057_l;
    reg node1058;
    reg node1059;
    reg node1060_r;
    reg node1060_l;
    reg node1061_r;
    reg node1061_l;
    reg node1062_r;
    reg node1062_l;
    reg node1063_r;
    reg node1063_l;
    reg node1064_r;
    reg node1064_l;
    reg node1065;
    reg node1066;
    reg node1067_r;
    reg node1067_l;
    reg node1068;
    reg node1069;
    reg node1070_r;
    reg node1070_l;
    reg node1071_r;
    reg node1071_l;
    reg node1072;
    reg node1073;
    reg node1074_r;
    reg node1074_l;
    reg node1075;
    reg node1076;
    reg node1077_r;
    reg node1077_l;
    reg node1078_r;
    reg node1078_l;
    reg node1079_r;
    reg node1079_l;
    reg node1080;
    reg node1081;
    reg node1082_r;
    reg node1082_l;
    reg node1083;
    reg node1084;
    reg node1085_r;
    reg node1085_l;
    reg node1086;
    reg node1087_r;
    reg node1087_l;
    reg node1088;
    reg node1089;
    reg node1090_r;
    reg node1090_l;
    reg node1091_r;
    reg node1091_l;
    reg node1092_r;
    reg node1092_l;
    reg node1093_r;
    reg node1093_l;
    reg node1094;
    reg node1095;
    reg node1096_r;
    reg node1096_l;
    reg node1097;
    reg node1098;
    reg node1099_r;
    reg node1099_l;
    reg node1100_r;
    reg node1100_l;
    reg node1101;
    reg node1102;
    reg node1103_r;
    reg node1103_l;
    reg node1104;
    reg node1105;
    reg node1106_r;
    reg node1106_l;
    reg node1107_r;
    reg node1107_l;
    reg node1108_r;
    reg node1108_l;
    reg node1109;
    reg node1110;
    reg node1111_r;
    reg node1111_l;
    reg node1112;
    reg node1113;
    reg node1114_r;
    reg node1114_l;
    reg node1115;
    reg node1116_r;
    reg node1116_l;
    reg node1117;
    reg node1118;
    reg node1119_r;
    reg node1119_l;
    reg node1120_r;
    reg node1120_l;
    reg node1121_r;
    reg node1121_l;
    reg node1122_r;
    reg node1122_l;
    reg node1123_r;
    reg node1123_l;
    reg node1124_r;
    reg node1124_l;
    reg node1125_r;
    reg node1125_l;
    reg node1126;
    reg node1127;
    reg node1128_r;
    reg node1128_l;
    reg node1129;
    reg node1130;
    reg node1131_r;
    reg node1131_l;
    reg node1132_r;
    reg node1132_l;
    reg node1133;
    reg node1134;
    reg node1135_r;
    reg node1135_l;
    reg node1136;
    reg node1137;
    reg node1138_r;
    reg node1138_l;
    reg node1139_r;
    reg node1139_l;
    reg node1140_r;
    reg node1140_l;
    reg node1141;
    reg node1142;
    reg node1143_r;
    reg node1143_l;
    reg node1144;
    reg node1145;
    reg node1146_r;
    reg node1146_l;
    reg node1147;
    reg node1148_r;
    reg node1148_l;
    reg node1149;
    reg node1150;
    reg node1151_r;
    reg node1151_l;
    reg node1152_r;
    reg node1152_l;
    reg node1153_r;
    reg node1153_l;
    reg node1154_r;
    reg node1154_l;
    reg node1155;
    reg node1156;
    reg node1157_r;
    reg node1157_l;
    reg node1158;
    reg node1159;
    reg node1160_r;
    reg node1160_l;
    reg node1161_r;
    reg node1161_l;
    reg node1162;
    reg node1163;
    reg node1164;
    reg node1165_r;
    reg node1165_l;
    reg node1166_r;
    reg node1166_l;
    reg node1167_r;
    reg node1167_l;
    reg node1168;
    reg node1169;
    reg node1170_r;
    reg node1170_l;
    reg node1171;
    reg node1172;
    reg node1173_r;
    reg node1173_l;
    reg node1174;
    reg node1175_r;
    reg node1175_l;
    reg node1176;
    reg node1177;
    reg node1178_r;
    reg node1178_l;
    reg node1179_r;
    reg node1179_l;
    reg node1180_r;
    reg node1180_l;
    reg node1181_r;
    reg node1181_l;
    reg node1182_r;
    reg node1182_l;
    reg node1183;
    reg node1184;
    reg node1185_r;
    reg node1185_l;
    reg node1186;
    reg node1187;
    reg node1188_r;
    reg node1188_l;
    reg node1189_r;
    reg node1189_l;
    reg node1190;
    reg node1191;
    reg node1192_r;
    reg node1192_l;
    reg node1193;
    reg node1194;
    reg node1195_r;
    reg node1195_l;
    reg node1196_r;
    reg node1196_l;
    reg node1197_r;
    reg node1197_l;
    reg node1198;
    reg node1199;
    reg node1200_r;
    reg node1200_l;
    reg node1201;
    reg node1202;
    reg node1203_r;
    reg node1203_l;
    reg node1204_r;
    reg node1204_l;
    reg node1205;
    reg node1206;
    reg node1207_r;
    reg node1207_l;
    reg node1208;
    reg node1209;
    reg node1210_r;
    reg node1210_l;
    reg node1211_r;
    reg node1211_l;
    reg node1212_r;
    reg node1212_l;
    reg node1213_r;
    reg node1213_l;
    reg node1214;
    reg node1215;
    reg node1216_r;
    reg node1216_l;
    reg node1217;
    reg node1218;
    reg node1219_r;
    reg node1219_l;
    reg node1220_r;
    reg node1220_l;
    reg node1221;
    reg node1222;
    reg node1223_r;
    reg node1223_l;
    reg node1224;
    reg node1225;
    reg node1226_r;
    reg node1226_l;
    reg node1227_r;
    reg node1227_l;
    reg node1228_r;
    reg node1228_l;
    reg node1229;
    reg node1230;
    reg node1231_r;
    reg node1231_l;
    reg node1232;
    reg node1233;
    reg node1234_r;
    reg node1234_l;
    reg node1235_r;
    reg node1235_l;
    reg node1236;
    reg node1237;
    reg node1238_r;
    reg node1238_l;
    reg node1239;
    reg node1240;
    reg node1241_r;
    reg node1241_l;
    reg node1242_r;
    reg node1242_l;
    reg node1243_r;
    reg node1243_l;
    reg node1244_r;
    reg node1244_l;
    reg node1245_r;
    reg node1245_l;
    reg node1246_r;
    reg node1246_l;
    reg node1247;
    reg node1248;
    reg node1249_r;
    reg node1249_l;
    reg node1250;
    reg node1251;
    reg node1252_r;
    reg node1252_l;
    reg node1253_r;
    reg node1253_l;
    reg node1254;
    reg node1255;
    reg node1256_r;
    reg node1256_l;
    reg node1257;
    reg node1258;
    reg node1259_r;
    reg node1259_l;
    reg node1260_r;
    reg node1260_l;
    reg node1261;
    reg node1262_r;
    reg node1262_l;
    reg node1263;
    reg node1264;
    reg node1265;
    reg node1266_r;
    reg node1266_l;
    reg node1267_r;
    reg node1267_l;
    reg node1268_r;
    reg node1268_l;
    reg node1269_r;
    reg node1269_l;
    reg node1270;
    reg node1271;
    reg node1272_r;
    reg node1272_l;
    reg node1273;
    reg node1274;
    reg node1275_r;
    reg node1275_l;
    reg node1276_r;
    reg node1276_l;
    reg node1277;
    reg node1278;
    reg node1279;
    reg node1280_r;
    reg node1280_l;
    reg node1281_r;
    reg node1281_l;
    reg node1282;
    reg node1283_r;
    reg node1283_l;
    reg node1284;
    reg node1285;
    reg node1286_r;
    reg node1286_l;
    reg node1287_r;
    reg node1287_l;
    reg node1288;
    reg node1289;
    reg node1290_r;
    reg node1290_l;
    reg node1291;
    reg node1292;
    reg node1293_r;
    reg node1293_l;
    reg node1294_r;
    reg node1294_l;
    reg node1295_r;
    reg node1295_l;
    reg node1296_r;
    reg node1296_l;
    reg node1297_r;
    reg node1297_l;
    reg node1298;
    reg node1299;
    reg node1300_r;
    reg node1300_l;
    reg node1301;
    reg node1302;
    reg node1303_r;
    reg node1303_l;
    reg node1304_r;
    reg node1304_l;
    reg node1305;
    reg node1306;
    reg node1307_r;
    reg node1307_l;
    reg node1308;
    reg node1309;
    reg node1310_r;
    reg node1310_l;
    reg node1311_r;
    reg node1311_l;
    reg node1312;
    reg node1313_r;
    reg node1313_l;
    reg node1314;
    reg node1315;
    reg node1316_r;
    reg node1316_l;
    reg node1317_r;
    reg node1317_l;
    reg node1318;
    reg node1319;
    reg node1320_r;
    reg node1320_l;
    reg node1321;
    reg node1322;
    reg node1323_r;
    reg node1323_l;
    reg node1324_r;
    reg node1324_l;
    reg node1325_r;
    reg node1325_l;
    reg node1326_r;
    reg node1326_l;
    reg node1327;
    reg node1328;
    reg node1329_r;
    reg node1329_l;
    reg node1330;
    reg node1331;
    reg node1332_r;
    reg node1332_l;
    reg node1333;
    reg node1334;
    reg node1335_r;
    reg node1335_l;
    reg node1336_r;
    reg node1336_l;
    reg node1337_r;
    reg node1337_l;
    reg node1338;
    reg node1339;
    reg node1340_r;
    reg node1340_l;
    reg node1341;
    reg node1342;
    reg node1343_r;
    reg node1343_l;
    reg node1344_r;
    reg node1344_l;
    reg node1345;
    reg node1346;
    reg node1347_r;
    reg node1347_l;
    reg node1348;
    reg node1349;
    reg node1350_r;
    reg node1350_l;
    reg node1351_r;
    reg node1351_l;
    reg node1352_r;
    reg node1352_l;
    reg node1353_r;
    reg node1353_l;
    reg node1354_r;
    reg node1354_l;
    reg node1355_r;
    reg node1355_l;
    reg node1356_r;
    reg node1356_l;
    reg node1357_r;
    reg node1357_l;
    reg node1358;
    reg node1359;
    reg node1360_r;
    reg node1360_l;
    reg node1361;
    reg node1362;
    reg node1363_r;
    reg node1363_l;
    reg node1364_r;
    reg node1364_l;
    reg node1365;
    reg node1366;
    reg node1367;
    reg node1368;
    reg node1369_r;
    reg node1369_l;
    reg node1370_r;
    reg node1370_l;
    reg node1371_r;
    reg node1371_l;
    reg node1372_r;
    reg node1372_l;
    reg node1373;
    reg node1374;
    reg node1375;
    reg node1376_r;
    reg node1376_l;
    reg node1377;
    reg node1378_r;
    reg node1378_l;
    reg node1379;
    reg node1380;
    reg node1381_r;
    reg node1381_l;
    reg node1382_r;
    reg node1382_l;
    reg node1383_r;
    reg node1383_l;
    reg node1384;
    reg node1385;
    reg node1386_r;
    reg node1386_l;
    reg node1387;
    reg node1388;
    reg node1389;
    reg node1390_r;
    reg node1390_l;
    reg node1391_r;
    reg node1391_l;
    reg node1392_r;
    reg node1392_l;
    reg node1393_r;
    reg node1393_l;
    reg node1394_r;
    reg node1394_l;
    reg node1395;
    reg node1396;
    reg node1397;
    reg node1398;
    reg node1399_r;
    reg node1399_l;
    reg node1400;
    reg node1401;
    reg node1402_r;
    reg node1402_l;
    reg node1403_r;
    reg node1403_l;
    reg node1404;
    reg node1405_r;
    reg node1405_l;
    reg node1406_r;
    reg node1406_l;
    reg node1407;
    reg node1408;
    reg node1409;
    reg node1410_r;
    reg node1410_l;
    reg node1411_r;
    reg node1411_l;
    reg node1412;
    reg node1413_r;
    reg node1413_l;
    reg node1414;
    reg node1415;
    reg node1416_r;
    reg node1416_l;
    reg node1417_r;
    reg node1417_l;
    reg node1418;
    reg node1419;
    reg node1420;
    reg node1421_r;
    reg node1421_l;
    reg node1422_r;
    reg node1422_l;
    reg node1423_r;
    reg node1423_l;
    reg node1424_r;
    reg node1424_l;
    reg node1425_r;
    reg node1425_l;
    reg node1426_r;
    reg node1426_l;
    reg node1427;
    reg node1428;
    reg node1429_r;
    reg node1429_l;
    reg node1430;
    reg node1431;
    reg node1432_r;
    reg node1432_l;
    reg node1433_r;
    reg node1433_l;
    reg node1434;
    reg node1435;
    reg node1436;
    reg node1437_r;
    reg node1437_l;
    reg node1438_r;
    reg node1438_l;
    reg node1439;
    reg node1440_r;
    reg node1440_l;
    reg node1441;
    reg node1442;
    reg node1443_r;
    reg node1443_l;
    reg node1444;
    reg node1445_r;
    reg node1445_l;
    reg node1446;
    reg node1447;
    reg node1448_r;
    reg node1448_l;
    reg node1449_r;
    reg node1449_l;
    reg node1450_r;
    reg node1450_l;
    reg node1451_r;
    reg node1451_l;
    reg node1452;
    reg node1453;
    reg node1454;
    reg node1455_r;
    reg node1455_l;
    reg node1456_r;
    reg node1456_l;
    reg node1457;
    reg node1458;
    reg node1459;
    reg node1460_r;
    reg node1460_l;
    reg node1461_r;
    reg node1461_l;
    reg node1462_r;
    reg node1462_l;
    reg node1463;
    reg node1464;
    reg node1465_r;
    reg node1465_l;
    reg node1466;
    reg node1467;
    reg node1468_r;
    reg node1468_l;
    reg node1469_r;
    reg node1469_l;
    reg node1470;
    reg node1471;
    reg node1472_r;
    reg node1472_l;
    reg node1473;
    reg node1474;
    reg node1475;
    reg node1476_r;
    reg node1476_l;
    reg node1477_r;
    reg node1477_l;
    reg node1478_r;
    reg node1478_l;
    reg node1479_r;
    reg node1479_l;
    reg node1480_r;
    reg node1480_l;
    reg node1481;
    reg node1482;
    reg node1483_r;
    reg node1483_l;
    reg node1484;
    reg node1485;
    reg node1486_r;
    reg node1486_l;
    reg node1487_r;
    reg node1487_l;
    reg node1488_r;
    reg node1488_l;
    reg node1489;
    reg node1490;
    reg node1491_r;
    reg node1491_l;
    reg node1492;
    reg node1493;
    reg node1494_r;
    reg node1494_l;
    reg node1495_r;
    reg node1495_l;
    reg node1496_r;
    reg node1496_l;
    reg node1497;
    reg node1498;
    reg node1499_r;
    reg node1499_l;
    reg node1500;
    reg node1501;
    reg node1502_r;
    reg node1502_l;
    reg node1503;
    reg node1504_r;
    reg node1504_l;
    reg node1505;
    reg node1506;
    reg node1507_r;
    reg node1507_l;
    reg node1508_r;
    reg node1508_l;
    reg node1509_r;
    reg node1509_l;
    reg node1510_r;
    reg node1510_l;
    reg node1511_r;
    reg node1511_l;
    reg node1512;
    reg node1513;
    reg node1514;
    reg node1515;
    reg node1516_r;
    reg node1516_l;
    reg node1517;
    reg node1518;
    reg node1519_r;
    reg node1519_l;
    reg node1520_r;
    reg node1520_l;
    reg node1521;
    reg node1522_r;
    reg node1522_l;
    reg node1523;
    reg node1524_r;
    reg node1524_l;
    reg node1525;
    reg node1526;
    reg node1527_r;
    reg node1527_l;
    reg node1528;
    reg node1529_r;
    reg node1529_l;
    reg node1530;
    reg node1531;
    reg node1532_r;
    reg node1532_l;
    reg node1533_r;
    reg node1533_l;
    reg node1534_r;
    reg node1534_l;
    reg node1535_r;
    reg node1535_l;
    reg node1536_r;
    reg node1536_l;
    reg node1537_r;
    reg node1537_l;
    reg node1538;
    reg node1539;
    reg node1540_r;
    reg node1540_l;
    reg node1541;
    reg node1542;
    reg node1543;
    reg node1544_r;
    reg node1544_l;
    reg node1545_r;
    reg node1545_l;
    reg node1546_r;
    reg node1546_l;
    reg node1547;
    reg node1548;
    reg node1549;
    reg node1550;
    reg node1551_r;
    reg node1551_l;
    reg node1552_r;
    reg node1552_l;
    reg node1553_r;
    reg node1553_l;
    reg node1554_r;
    reg node1554_l;
    reg node1555;
    reg node1556;
    reg node1557;
    reg node1558_r;
    reg node1558_l;
    reg node1559;
    reg node1560;
    reg node1561_r;
    reg node1561_l;
    reg node1562_r;
    reg node1562_l;
    reg node1563;
    reg node1564;
    reg node1565_r;
    reg node1565_l;
    reg node1566_r;
    reg node1566_l;
    reg node1567;
    reg node1568;
    reg node1569;
    reg node1570_r;
    reg node1570_l;
    reg node1571_r;
    reg node1571_l;
    reg node1572_r;
    reg node1572_l;
    reg node1573_r;
    reg node1573_l;
    reg node1574_r;
    reg node1574_l;
    reg node1575;
    reg node1576;
    reg node1577_r;
    reg node1577_l;
    reg node1578;
    reg node1579;
    reg node1580_r;
    reg node1580_l;
    reg node1581_r;
    reg node1581_l;
    reg node1582;
    reg node1583;
    reg node1584;
    reg node1585_r;
    reg node1585_l;
    reg node1586_r;
    reg node1586_l;
    reg node1587;
    reg node1588;
    reg node1589;
    reg node1590_r;
    reg node1590_l;
    reg node1591_r;
    reg node1591_l;
    reg node1592_r;
    reg node1592_l;
    reg node1593_r;
    reg node1593_l;
    reg node1594;
    reg node1595;
    reg node1596_r;
    reg node1596_l;
    reg node1597;
    reg node1598;
    reg node1599;
    reg node1600_r;
    reg node1600_l;
    reg node1601_r;
    reg node1601_l;
    reg node1602;
    reg node1603_r;
    reg node1603_l;
    reg node1604;
    reg node1605;
    reg node1606_r;
    reg node1606_l;
    reg node1607_r;
    reg node1607_l;
    reg node1608;
    reg node1609;
    reg node1610_r;
    reg node1610_l;
    reg node1611;
    reg node1612;
    reg result0;
    reg result1;
    reg result2;
    reg result3;
    reg result4;
    reg result5;
    reg result6;
    reg result7;
    reg result8;
    reg result9;

    begin
      node0_r = pixel[568];
      node0_l = ~pixel[568];
      node1_r = node0_l & pixel[430];
      node1_l = node0_l & ~pixel[430];
      node2_r = node1_l & pixel[378];
      node2_l = node1_l & ~pixel[378];
      node3_r = node2_l & pixel[487];
      node3_l = node2_l & ~pixel[487];
      node4_r = node3_l & pixel[566];
      node4_l = node3_l & ~pixel[566];
      node5_r = node4_l & pixel[182];
      node5_l = node4_l & ~pixel[182];
      node6_r = node5_l & pixel[95];
      node6_l = node5_l & ~pixel[95];
      node7_r = node6_l & pixel[158];
      node7_l = node6_l & ~pixel[158];
      node8_r = node7_l & pixel[512];
      node8_l = node7_l & ~pixel[512];
      node9_r = node8_l & pixel[431];
      node9_l = node8_l & ~pixel[431];
      node10 = node9_l;
      node11 = node9_r;
      node12_r = node8_r & pixel[98];
      node12_l = node8_r & ~pixel[98];
      node13 = node12_l;
      node14 = node12_r;
      node15_r = node7_r & pixel[326];
      node15_l = node7_r & ~pixel[326];
      node16_r = node15_l & pixel[330];
      node16_l = node15_l & ~pixel[330];
      node17 = node16_l;
      node18 = node16_r;
      node19_r = node15_r & pixel[599];
      node19_l = node15_r & ~pixel[599];
      node20 = node19_l;
      node21 = node19_r;
      node22_r = node6_r & pixel[498];
      node22_l = node6_r & ~pixel[498];
      node23_r = node22_l & pixel[629];
      node23_l = node22_l & ~pixel[629];
      node24 = node23_l;
      node25 = node23_r;
      node26 = node22_r;
      node27_r = node5_r & pixel[660];
      node27_l = node5_r & ~pixel[660];
      node28_r = node27_l & pixel[633];
      node28_l = node27_l & ~pixel[633];
      node29_r = node28_l & pixel[269];
      node29_l = node28_l & ~pixel[269];
      node30_r = node29_l & pixel[709];
      node30_l = node29_l & ~pixel[709];
      node31 = node30_l;
      node32 = node30_r;
      node33_r = node29_r & pixel[299];
      node33_l = node29_r & ~pixel[299];
      node34 = node33_l;
      node35 = node33_r;
      node36_r = node28_r & pixel[626];
      node36_l = node28_r & ~pixel[626];
      node37_r = node36_l & pixel[437];
      node37_l = node36_l & ~pixel[437];
      node38 = node37_l;
      node39 = node37_r;
      node40_r = node36_r & pixel[498];
      node40_l = node36_r & ~pixel[498];
      node41 = node40_l;
      node42 = node40_r;
      node43_r = node27_r & pixel[513];
      node43_l = node27_r & ~pixel[513];
      node44_r = node43_l & pixel[404];
      node44_l = node43_l & ~pixel[404];
      node45_r = node44_l & pixel[345];
      node45_l = node44_l & ~pixel[345];
      node46 = node45_l;
      node47 = node45_r;
      node48_r = node44_r & pixel[517];
      node48_l = node44_r & ~pixel[517];
      node49 = node48_l;
      node50 = node48_r;
      node51_r = node43_r & pixel[635];
      node51_l = node43_r & ~pixel[635];
      node52_r = node51_l & pixel[259];
      node52_l = node51_l & ~pixel[259];
      node53 = node52_l;
      node54 = node52_r;
      node55_r = node51_r & pixel[129];
      node55_l = node51_r & ~pixel[129];
      node56 = node55_l;
      node57 = node55_r;
      node58_r = node4_r & pixel[178];
      node58_l = node4_r & ~pixel[178];
      node59_r = node58_l & pixel[426];
      node59_l = node58_l & ~pixel[426];
      node60_r = node59_l & pixel[399];
      node60_l = node59_l & ~pixel[399];
      node61_r = node60_l & pixel[126];
      node61_l = node60_l & ~pixel[126];
      node62_r = node61_l & pixel[264];
      node62_l = node61_l & ~pixel[264];
      node63 = node62_l;
      node64 = node62_r;
      node65_r = node61_r & pixel[133];
      node65_l = node61_r & ~pixel[133];
      node66 = node65_l;
      node67 = node65_r;
      node68_r = node60_r & pixel[205];
      node68_l = node60_r & ~pixel[205];
      node69 = node68_l;
      node70 = node68_r;
      node71_r = node59_r & pixel[715];
      node71_l = node59_r & ~pixel[715];
      node72_r = node71_l & pixel[323];
      node72_l = node71_l & ~pixel[323];
      node73 = node72_l;
      node74_r = node72_r & pixel[163];
      node74_l = node72_r & ~pixel[163];
      node75 = node74_l;
      node76 = node74_r;
      node77_r = node71_r & pixel[443];
      node77_l = node71_r & ~pixel[443];
      node78 = node77_l;
      node79 = node77_r;
      node80_r = node58_r & pixel[302];
      node80_l = node58_r & ~pixel[302];
      node81_r = node80_l & pixel[342];
      node81_l = node80_l & ~pixel[342];
      node82_r = node81_l & pixel[220];
      node82_l = node81_l & ~pixel[220];
      node83_r = node82_l & pixel[428];
      node83_l = node82_l & ~pixel[428];
      node84 = node83_l;
      node85 = node83_r;
      node86 = node82_r;
      node87_r = node81_r & pixel[341];
      node87_l = node81_r & ~pixel[341];
      node88_r = node87_l & pixel[243];
      node88_l = node87_l & ~pixel[243];
      node89 = node88_l;
      node90 = node88_r;
      node91 = node87_r;
      node92_r = node80_r & pixel[228];
      node92_l = node80_r & ~pixel[228];
      node93 = node92_l;
      node94 = node92_r;
      node95_r = node3_r & pixel[626];
      node95_l = node3_r & ~pixel[626];
      node96_r = node95_l & pixel[455];
      node96_l = node95_l & ~pixel[455];
      node97_r = node96_l & pixel[353];
      node97_l = node96_l & ~pixel[353];
      node98_r = node97_l & pixel[377];
      node98_l = node97_l & ~pixel[377];
      node99_r = node98_l & pixel[98];
      node99_l = node98_l & ~pixel[98];
      node100_r = node99_l & pixel[191];
      node100_l = node99_l & ~pixel[191];
      node101 = node100_l;
      node102 = node100_r;
      node103 = node99_r;
      node104_r = node98_r & pixel[686];
      node104_l = node98_r & ~pixel[686];
      node105_r = node104_l & pixel[179];
      node105_l = node104_l & ~pixel[179];
      node106 = node105_l;
      node107 = node105_r;
      node108 = node104_r;
      node109_r = node97_r & pixel[429];
      node109_l = node97_r & ~pixel[429];
      node110_r = node109_l & pixel[493];
      node110_l = node109_l & ~pixel[493];
      node111_r = node110_l & pixel[629];
      node111_l = node110_l & ~pixel[629];
      node112 = node111_l;
      node113 = node111_r;
      node114_r = node110_r & pixel[374];
      node114_l = node110_r & ~pixel[374];
      node115 = node114_l;
      node116 = node114_r;
      node117_r = node109_r & pixel[357];
      node117_l = node109_r & ~pixel[357];
      node118_r = node117_l & pixel[496];
      node118_l = node117_l & ~pixel[496];
      node119 = node118_l;
      node120 = node118_r;
      node121 = node117_r;
      node122_r = node96_r & pixel[241];
      node122_l = node96_r & ~pixel[241];
      node123_r = node122_l & pixel[554];
      node123_l = node122_l & ~pixel[554];
      node124_r = node123_l & pixel[184];
      node124_l = node123_l & ~pixel[184];
      node125_r = node124_l & pixel[153];
      node125_l = node124_l & ~pixel[153];
      node126 = node125_l;
      node127 = node125_r;
      node128_r = node124_r & pixel[212];
      node128_l = node124_r & ~pixel[212];
      node129 = node128_l;
      node130 = node128_r;
      node131_r = node123_r & pixel[216];
      node131_l = node123_r & ~pixel[216];
      node132_r = node131_l & pixel[574];
      node132_l = node131_l & ~pixel[574];
      node133 = node132_l;
      node134 = node132_r;
      node135_r = node131_r & pixel[551];
      node135_l = node131_r & ~pixel[551];
      node136 = node135_l;
      node137 = node135_r;
      node138_r = node122_r & pixel[209];
      node138_l = node122_r & ~pixel[209];
      node139_r = node138_l & pixel[523];
      node139_l = node138_l & ~pixel[523];
      node140_r = node139_l & pixel[741];
      node140_l = node139_l & ~pixel[741];
      node141 = node140_l;
      node142 = node140_r;
      node143_r = node139_r & pixel[485];
      node143_l = node139_r & ~pixel[485];
      node144 = node143_l;
      node145 = node143_r;
      node146_r = node138_r & pixel[441];
      node146_l = node138_r & ~pixel[441];
      node147_r = node146_l & pixel[249];
      node147_l = node146_l & ~pixel[249];
      node148 = node147_l;
      node149 = node147_r;
      node150_r = node146_r & pixel[347];
      node150_l = node146_r & ~pixel[347];
      node151 = node150_l;
      node152 = node150_r;
      node153_r = node95_r & pixel[374];
      node153_l = node95_r & ~pixel[374];
      node154_r = node153_l & pixel[376];
      node154_l = node153_l & ~pixel[376];
      node155_r = node154_l & pixel[680];
      node155_l = node154_l & ~pixel[680];
      node156_r = node155_l & pixel[399];
      node156_l = node155_l & ~pixel[399];
      node157_r = node156_l & pixel[373];
      node157_l = node156_l & ~pixel[373];
      node158 = node157_l;
      node159 = node157_r;
      node160_r = node156_r & pixel[267];
      node160_l = node156_r & ~pixel[267];
      node161 = node160_l;
      node162 = node160_r;
      node163_r = node155_r & pixel[598];
      node163_l = node155_r & ~pixel[598];
      node164_r = node163_l & pixel[186];
      node164_l = node163_l & ~pixel[186];
      node165 = node164_l;
      node166 = node164_r;
      node167_r = node163_r & pixel[464];
      node167_l = node163_r & ~pixel[464];
      node168 = node167_l;
      node169 = node167_r;
      node170_r = node154_r & pixel[522];
      node170_l = node154_r & ~pixel[522];
      node171_r = node170_l & pixel[96];
      node171_l = node170_l & ~pixel[96];
      node172_r = node171_l & pixel[681];
      node172_l = node171_l & ~pixel[681];
      node173 = node172_l;
      node174 = node172_r;
      node175 = node171_r;
      node176_r = node170_r & pixel[323];
      node176_l = node170_r & ~pixel[323];
      node177 = node176_l;
      node178 = node176_r;
      node179_r = node153_r & pixel[405];
      node179_l = node153_r & ~pixel[405];
      node180_r = node179_l & pixel[240];
      node180_l = node179_l & ~pixel[240];
      node181_r = node180_l & pixel[601];
      node181_l = node180_l & ~pixel[601];
      node182_r = node181_l & pixel[372];
      node182_l = node181_l & ~pixel[372];
      node183 = node182_l;
      node184 = node182_r;
      node185 = node181_r;
      node186_r = node180_r & pixel[435];
      node186_l = node180_r & ~pixel[435];
      node187 = node186_l;
      node188_r = node186_r & pixel[272];
      node188_l = node186_r & ~pixel[272];
      node189 = node188_l;
      node190 = node188_r;
      node191_r = node179_r & pixel[651];
      node191_l = node179_r & ~pixel[651];
      node192_r = node191_l & pixel[354];
      node192_l = node191_l & ~pixel[354];
      node193_r = node192_l & pixel[570];
      node193_l = node192_l & ~pixel[570];
      node194 = node193_l;
      node195 = node193_r;
      node196_r = node192_r & pixel[293];
      node196_l = node192_r & ~pixel[293];
      node197 = node196_l;
      node198 = node196_r;
      node199_r = node191_r & pixel[654];
      node199_l = node191_r & ~pixel[654];
      node200 = node199_l;
      node201_r = node199_r & pixel[571];
      node201_l = node199_r & ~pixel[571];
      node202 = node201_l;
      node203 = node201_r;
      node204_r = node2_r & pixel[354];
      node204_l = node2_r & ~pixel[354];
      node205_r = node204_l & pixel[437];
      node205_l = node204_l & ~pixel[437];
      node206_r = node205_l & pixel[522];
      node206_l = node205_l & ~pixel[522];
      node207_r = node206_l & pixel[325];
      node207_l = node206_l & ~pixel[325];
      node208_r = node207_l & pixel[191];
      node208_l = node207_l & ~pixel[191];
      node209_r = node208_l & pixel[290];
      node209_l = node208_l & ~pixel[290];
      node210_r = node209_l & pixel[580];
      node210_l = node209_l & ~pixel[580];
      node211 = node210_l;
      node212 = node210_r;
      node213_r = node209_r & pixel[681];
      node213_l = node209_r & ~pixel[681];
      node214 = node213_l;
      node215 = node213_r;
      node216_r = node208_r & pixel[217];
      node216_l = node208_r & ~pixel[217];
      node217_r = node216_l & pixel[439];
      node217_l = node216_l & ~pixel[439];
      node218 = node217_l;
      node219 = node217_r;
      node220 = node216_r;
      node221_r = node207_r & pixel[578];
      node221_l = node207_r & ~pixel[578];
      node222_r = node221_l & pixel[630];
      node222_l = node221_l & ~pixel[630];
      node223_r = node222_l & pixel[210];
      node223_l = node222_l & ~pixel[210];
      node224 = node223_l;
      node225 = node223_r;
      node226_r = node222_r & pixel[266];
      node226_l = node222_r & ~pixel[266];
      node227 = node226_l;
      node228 = node226_r;
      node229_r = node221_r & pixel[376];
      node229_l = node221_r & ~pixel[376];
      node230_r = node229_l & pixel[456];
      node230_l = node229_l & ~pixel[456];
      node231 = node230_l;
      node232 = node230_r;
      node233_r = node229_r & pixel[579];
      node233_l = node229_r & ~pixel[579];
      node234 = node233_l;
      node235 = node233_r;
      node236_r = node206_r & pixel[318];
      node236_l = node206_r & ~pixel[318];
      node237_r = node236_l & pixel[526];
      node237_l = node236_l & ~pixel[526];
      node238_r = node237_l & pixel[465];
      node238_l = node237_l & ~pixel[465];
      node239_r = node238_l & pixel[293];
      node239_l = node238_l & ~pixel[293];
      node240 = node239_l;
      node241 = node239_r;
      node242_r = node238_r & pixel[685];
      node242_l = node238_r & ~pixel[685];
      node243 = node242_l;
      node244 = node242_r;
      node245_r = node237_r & pixel[442];
      node245_l = node237_r & ~pixel[442];
      node246_r = node245_l & pixel[331];
      node246_l = node245_l & ~pixel[331];
      node247 = node246_l;
      node248 = node246_r;
      node249_r = node245_r & pixel[259];
      node249_l = node245_r & ~pixel[259];
      node250 = node249_l;
      node251 = node249_r;
      node252_r = node236_r & pixel[496];
      node252_l = node236_r & ~pixel[496];
      node253_r = node252_l & pixel[488];
      node253_l = node252_l & ~pixel[488];
      node254_r = node253_l & pixel[158];
      node254_l = node253_l & ~pixel[158];
      node255 = node254_l;
      node256 = node254_r;
      node257_r = node253_r & pixel[383];
      node257_l = node253_r & ~pixel[383];
      node258 = node257_l;
      node259 = node257_r;
      node260_r = node252_r & pixel[472];
      node260_l = node252_r & ~pixel[472];
      node261_r = node260_l & pixel[600];
      node261_l = node260_l & ~pixel[600];
      node262 = node261_l;
      node263 = node261_r;
      node264 = node260_r;
      node265_r = node205_r & pixel[151];
      node265_l = node205_r & ~pixel[151];
      node266_r = node265_l & pixel[296];
      node266_l = node265_l & ~pixel[296];
      node267_r = node266_l & pixel[102];
      node267_l = node266_l & ~pixel[102];
      node268_r = node267_l & pixel[262];
      node268_l = node267_l & ~pixel[262];
      node269_r = node268_l & pixel[263];
      node269_l = node268_l & ~pixel[263];
      node270 = node269_l;
      node271 = node269_r;
      node272_r = node268_r & pixel[295];
      node272_l = node268_r & ~pixel[295];
      node273 = node272_l;
      node274 = node272_r;
      node275 = node267_r;
      node276_r = node266_r & pixel[183];
      node276_l = node266_r & ~pixel[183];
      node277_r = node276_l & pixel[347];
      node277_l = node276_l & ~pixel[347];
      node278_r = node277_l & pixel[375];
      node278_l = node277_l & ~pixel[375];
      node279 = node278_l;
      node280 = node278_r;
      node281_r = node277_r & pixel[715];
      node281_l = node277_r & ~pixel[715];
      node282 = node281_l;
      node283 = node281_r;
      node284_r = node276_r & pixel[651];
      node284_l = node276_r & ~pixel[651];
      node285_r = node284_l & pixel[319];
      node285_l = node284_l & ~pixel[319];
      node286 = node285_l;
      node287 = node285_r;
      node288_r = node284_r & pixel[357];
      node288_l = node284_r & ~pixel[357];
      node289 = node288_l;
      node290 = node288_r;
      node291_r = node265_r & pixel[324];
      node291_l = node265_r & ~pixel[324];
      node292_r = node291_l & pixel[236];
      node292_l = node291_l & ~pixel[236];
      node293_r = node292_l & pixel[487];
      node293_l = node292_l & ~pixel[487];
      node294_r = node293_l & pixel[241];
      node294_l = node293_l & ~pixel[241];
      node295 = node294_l;
      node296 = node294_r;
      node297_r = node293_r & pixel[432];
      node297_l = node293_r & ~pixel[432];
      node298 = node297_l;
      node299 = node297_r;
      node300_r = node292_r & pixel[146];
      node300_l = node292_r & ~pixel[146];
      node301_r = node300_l & pixel[489];
      node301_l = node300_l & ~pixel[489];
      node302 = node301_l;
      node303 = node301_r;
      node304 = node300_r;
      node305_r = node291_r & pixel[622];
      node305_l = node291_r & ~pixel[622];
      node306_r = node305_l & pixel[625];
      node306_l = node305_l & ~pixel[625];
      node307_r = node306_l & pixel[460];
      node307_l = node306_l & ~pixel[460];
      node308 = node307_l;
      node309 = node307_r;
      node310_r = node306_r & pixel[545];
      node310_l = node306_r & ~pixel[545];
      node311 = node310_l;
      node312 = node310_r;
      node313_r = node305_r & pixel[190];
      node313_l = node305_r & ~pixel[190];
      node314_r = node313_l & pixel[621];
      node314_l = node313_l & ~pixel[621];
      node315 = node314_l;
      node316 = node314_r;
      node317_r = node313_r & pixel[293];
      node317_l = node313_r & ~pixel[293];
      node318 = node317_l;
      node319 = node317_r;
      node320_r = node204_r & pixel[595];
      node320_l = node204_r & ~pixel[595];
      node321_r = node320_l & pixel[460];
      node321_l = node320_l & ~pixel[460];
      node322_r = node321_l & pixel[184];
      node322_l = node321_l & ~pixel[184];
      node323_r = node322_l & pixel[485];
      node323_l = node322_l & ~pixel[485];
      node324_r = node323_l & pixel[240];
      node324_l = node323_l & ~pixel[240];
      node325_r = node324_l & pixel[287];
      node325_l = node324_l & ~pixel[287];
      node326 = node325_l;
      node327 = node325_r;
      node328_r = node324_r & pixel[376];
      node328_l = node324_r & ~pixel[376];
      node329 = node328_l;
      node330 = node328_r;
      node331_r = node323_r & pixel[122];
      node331_l = node323_r & ~pixel[122];
      node332_r = node331_l & pixel[293];
      node332_l = node331_l & ~pixel[293];
      node333 = node332_l;
      node334 = node332_r;
      node335 = node331_r;
      node336_r = node322_r & pixel[440];
      node336_l = node322_r & ~pixel[440];
      node337_r = node336_l & pixel[203];
      node337_l = node336_l & ~pixel[203];
      node338_r = node337_l & pixel[153];
      node338_l = node337_l & ~pixel[153];
      node339 = node338_l;
      node340 = node338_r;
      node341_r = node337_r & pixel[404];
      node341_l = node337_r & ~pixel[404];
      node342 = node341_l;
      node343 = node341_r;
      node344_r = node336_r & pixel[622];
      node344_l = node336_r & ~pixel[622];
      node345_r = node344_l & pixel[268];
      node345_l = node344_l & ~pixel[268];
      node346 = node345_l;
      node347 = node345_r;
      node348_r = node344_r & pixel[271];
      node348_l = node344_r & ~pixel[271];
      node349 = node348_l;
      node350 = node348_r;
      node351_r = node321_r & pixel[318];
      node351_l = node321_r & ~pixel[318];
      node352_r = node351_l & pixel[205];
      node352_l = node351_l & ~pixel[205];
      node353_r = node352_l & pixel[235];
      node353_l = node352_l & ~pixel[235];
      node354_r = node353_l & pixel[155];
      node354_l = node353_l & ~pixel[155];
      node355 = node354_l;
      node356 = node354_r;
      node357_r = node353_r & pixel[316];
      node357_l = node353_r & ~pixel[316];
      node358 = node357_l;
      node359 = node357_r;
      node360_r = node352_r & pixel[316];
      node360_l = node352_r & ~pixel[316];
      node361_r = node360_l & pixel[151];
      node361_l = node360_l & ~pixel[151];
      node362 = node361_l;
      node363 = node361_r;
      node364_r = node360_r & pixel[456];
      node364_l = node360_r & ~pixel[456];
      node365 = node364_l;
      node366 = node364_r;
      node367_r = node351_r & pixel[371];
      node367_l = node351_r & ~pixel[371];
      node368_r = node367_l & pixel[377];
      node368_l = node367_l & ~pixel[377];
      node369_r = node368_l & pixel[260];
      node369_l = node368_l & ~pixel[260];
      node370 = node369_l;
      node371 = node369_r;
      node372_r = node368_r & pixel[570];
      node372_l = node368_r & ~pixel[570];
      node373 = node372_l;
      node374 = node372_r;
      node375_r = node367_r & pixel[543];
      node375_l = node367_r & ~pixel[543];
      node376_r = node375_l & pixel[513];
      node376_l = node375_l & ~pixel[513];
      node377 = node376_l;
      node378 = node376_r;
      node379_r = node375_r & pixel[655];
      node379_l = node375_r & ~pixel[655];
      node380 = node379_l;
      node381 = node379_r;
      node382_r = node320_r & pixel[270];
      node382_l = node320_r & ~pixel[270];
      node383_r = node382_l & pixel[328];
      node383_l = node382_l & ~pixel[328];
      node384_r = node383_l & pixel[318];
      node384_l = node383_l & ~pixel[318];
      node385_r = node384_l & pixel[555];
      node385_l = node384_l & ~pixel[555];
      node386_r = node385_l & pixel[124];
      node386_l = node385_l & ~pixel[124];
      node387 = node386_l;
      node388 = node386_r;
      node389_r = node385_r & pixel[407];
      node389_l = node385_r & ~pixel[407];
      node390 = node389_l;
      node391 = node389_r;
      node392_r = node384_r & pixel[267];
      node392_l = node384_r & ~pixel[267];
      node393_r = node392_l & pixel[657];
      node393_l = node392_l & ~pixel[657];
      node394 = node393_l;
      node395 = node393_r;
      node396_r = node392_r & pixel[298];
      node396_l = node392_r & ~pixel[298];
      node397 = node396_l;
      node398 = node396_r;
      node399_r = node383_r & pixel[514];
      node399_l = node383_r & ~pixel[514];
      node400_r = node399_l & pixel[570];
      node400_l = node399_l & ~pixel[570];
      node401_r = node400_l & pixel[259];
      node401_l = node400_l & ~pixel[259];
      node402 = node401_l;
      node403 = node401_r;
      node404 = node400_r;
      node405 = node399_r;
      node406_r = node382_r & pixel[569];
      node406_l = node382_r & ~pixel[569];
      node407_r = node406_l & pixel[515];
      node407_l = node406_l & ~pixel[515];
      node408_r = node407_l & pixel[290];
      node408_l = node407_l & ~pixel[290];
      node409_r = node408_l & pixel[398];
      node409_l = node408_l & ~pixel[398];
      node410 = node409_l;
      node411 = node409_r;
      node412_r = node408_r & pixel[371];
      node412_l = node408_r & ~pixel[371];
      node413 = node412_l;
      node414 = node412_r;
      node415_r = node407_r & pixel[631];
      node415_l = node407_r & ~pixel[631];
      node416 = node415_l;
      node417 = node415_r;
      node418_r = node406_r & pixel[404];
      node418_l = node406_r & ~pixel[404];
      node419_r = node418_l & pixel[291];
      node419_l = node418_l & ~pixel[291];
      node420_r = node419_l & pixel[182];
      node420_l = node419_l & ~pixel[182];
      node421 = node420_l;
      node422 = node420_r;
      node423 = node419_r;
      node424_r = node418_r & pixel[246];
      node424_l = node418_r & ~pixel[246];
      node425 = node424_l;
      node426 = node424_r;
      node427_r = node1_r & pixel[542];
      node427_l = node1_r & ~pixel[542];
      node428_r = node427_l & pixel[317];
      node428_l = node427_l & ~pixel[317];
      node429_r = node428_l & pixel[463];
      node429_l = node428_l & ~pixel[463];
      node430_r = node429_l & pixel[179];
      node430_l = node429_l & ~pixel[179];
      node431_r = node430_l & pixel[320];
      node431_l = node430_l & ~pixel[320];
      node432_r = node431_l & pixel[237];
      node432_l = node431_l & ~pixel[237];
      node433_r = node432_l & pixel[624];
      node433_l = node432_l & ~pixel[624];
      node434_r = node433_l & pixel[258];
      node434_l = node433_l & ~pixel[258];
      node435 = node434_l;
      node436 = node434_r;
      node437_r = node433_r & pixel[406];
      node437_l = node433_r & ~pixel[406];
      node438 = node437_l;
      node439 = node437_r;
      node440_r = node432_r & pixel[185];
      node440_l = node432_r & ~pixel[185];
      node441_r = node440_l & pixel[517];
      node441_l = node440_l & ~pixel[517];
      node442 = node441_l;
      node443 = node441_r;
      node444_r = node440_r & pixel[608];
      node444_l = node440_r & ~pixel[608];
      node445 = node444_l;
      node446 = node444_r;
      node447_r = node431_r & pixel[655];
      node447_l = node431_r & ~pixel[655];
      node448_r = node447_l & pixel[578];
      node448_l = node447_l & ~pixel[578];
      node449_r = node448_l & pixel[627];
      node449_l = node448_l & ~pixel[627];
      node450 = node449_l;
      node451 = node449_r;
      node452_r = node448_r & pixel[689];
      node452_l = node448_r & ~pixel[689];
      node453 = node452_l;
      node454 = node452_r;
      node455_r = node447_r & pixel[442];
      node455_l = node447_r & ~pixel[442];
      node456_r = node455_l & pixel[385];
      node456_l = node455_l & ~pixel[385];
      node457 = node456_l;
      node458 = node456_r;
      node459_r = node455_r & pixel[623];
      node459_l = node455_r & ~pixel[623];
      node460 = node459_l;
      node461 = node459_r;
      node462_r = node430_r & pixel[342];
      node462_l = node430_r & ~pixel[342];
      node463_r = node462_l & pixel[210];
      node463_l = node462_l & ~pixel[210];
      node464_r = node463_l & pixel[241];
      node464_l = node463_l & ~pixel[241];
      node465_r = node464_l & pixel[545];
      node465_l = node464_l & ~pixel[545];
      node466 = node465_l;
      node467 = node465_r;
      node468_r = node464_r & pixel[482];
      node468_l = node464_r & ~pixel[482];
      node469 = node468_l;
      node470 = node468_r;
      node471_r = node463_r & pixel[325];
      node471_l = node463_r & ~pixel[325];
      node472_r = node471_l & pixel[217];
      node472_l = node471_l & ~pixel[217];
      node473 = node472_l;
      node474 = node472_r;
      node475_r = node471_r & pixel[511];
      node475_l = node471_r & ~pixel[511];
      node476 = node475_l;
      node477 = node475_r;
      node478_r = node462_r & pixel[186];
      node478_l = node462_r & ~pixel[186];
      node479_r = node478_l & pixel[414];
      node479_l = node478_l & ~pixel[414];
      node480_r = node479_l & pixel[181];
      node480_l = node479_l & ~pixel[181];
      node481 = node480_l;
      node482 = node480_r;
      node483_r = node479_r & pixel[398];
      node483_l = node479_r & ~pixel[398];
      node484 = node483_l;
      node485 = node483_r;
      node486_r = node478_r & pixel[298];
      node486_l = node478_r & ~pixel[298];
      node487_r = node486_l & pixel[628];
      node487_l = node486_l & ~pixel[628];
      node488 = node487_l;
      node489 = node487_r;
      node490_r = node486_r & pixel[182];
      node490_l = node486_r & ~pixel[182];
      node491 = node490_l;
      node492 = node490_r;
      node493_r = node429_r & pixel[624];
      node493_l = node429_r & ~pixel[624];
      node494_r = node493_l & pixel[179];
      node494_l = node493_l & ~pixel[179];
      node495_r = node494_l & pixel[456];
      node495_l = node494_l & ~pixel[456];
      node496_r = node495_l & pixel[494];
      node496_l = node495_l & ~pixel[494];
      node497_r = node496_l & pixel[711];
      node497_l = node496_l & ~pixel[711];
      node498 = node497_l;
      node499 = node497_r;
      node500_r = node496_r & pixel[232];
      node500_l = node496_r & ~pixel[232];
      node501 = node500_l;
      node502 = node500_r;
      node503_r = node495_r & pixel[235];
      node503_l = node495_r & ~pixel[235];
      node504_r = node503_l & pixel[467];
      node504_l = node503_l & ~pixel[467];
      node505 = node504_l;
      node506 = node504_r;
      node507_r = node503_r & pixel[342];
      node507_l = node503_r & ~pixel[342];
      node508 = node507_l;
      node509 = node507_r;
      node510_r = node494_r & pixel[314];
      node510_l = node494_r & ~pixel[314];
      node511_r = node510_l & pixel[295];
      node511_l = node510_l & ~pixel[295];
      node512_r = node511_l & pixel[210];
      node512_l = node511_l & ~pixel[210];
      node513 = node512_l;
      node514 = node512_r;
      node515_r = node511_r & pixel[545];
      node515_l = node511_r & ~pixel[545];
      node516 = node515_l;
      node517 = node515_r;
      node518_r = node510_r & pixel[411];
      node518_l = node510_r & ~pixel[411];
      node519_r = node518_l & pixel[551];
      node519_l = node518_l & ~pixel[551];
      node520 = node519_l;
      node521 = node519_r;
      node522_r = node518_r & pixel[267];
      node522_l = node518_r & ~pixel[267];
      node523 = node522_l;
      node524 = node522_r;
      node525_r = node493_r & pixel[379];
      node525_l = node493_r & ~pixel[379];
      node526_r = node525_l & pixel[375];
      node526_l = node525_l & ~pixel[375];
      node527_r = node526_l & pixel[510];
      node527_l = node526_l & ~pixel[510];
      node528_r = node527_l & pixel[412];
      node528_l = node527_l & ~pixel[412];
      node529 = node528_l;
      node530 = node528_r;
      node531 = node527_r;
      node532_r = node526_r & pixel[154];
      node532_l = node526_r & ~pixel[154];
      node533_r = node532_l & pixel[411];
      node533_l = node532_l & ~pixel[411];
      node534 = node533_l;
      node535 = node533_r;
      node536_r = node532_r & pixel[301];
      node536_l = node532_r & ~pixel[301];
      node537 = node536_l;
      node538 = node536_r;
      node539_r = node525_r & pixel[320];
      node539_l = node525_r & ~pixel[320];
      node540_r = node539_l & pixel[512];
      node540_l = node539_l & ~pixel[512];
      node541_r = node540_l & pixel[652];
      node541_l = node540_l & ~pixel[652];
      node542 = node541_l;
      node543 = node541_r;
      node544_r = node540_r & pixel[575];
      node544_l = node540_r & ~pixel[575];
      node545 = node544_l;
      node546 = node544_r;
      node547_r = node539_r & pixel[483];
      node547_l = node539_r & ~pixel[483];
      node548_r = node547_l & pixel[245];
      node548_l = node547_l & ~pixel[245];
      node549 = node548_l;
      node550 = node548_r;
      node551_r = node547_r & pixel[301];
      node551_l = node547_r & ~pixel[301];
      node552 = node551_l;
      node553 = node551_r;
      node554_r = node428_r & pixel[211];
      node554_l = node428_r & ~pixel[211];
      node555_r = node554_l & pixel[96];
      node555_l = node554_l & ~pixel[96];
      node556_r = node555_l & pixel[322];
      node556_l = node555_l & ~pixel[322];
      node557_r = node556_l & pixel[237];
      node557_l = node556_l & ~pixel[237];
      node558_r = node557_l & pixel[651];
      node558_l = node557_l & ~pixel[651];
      node559_r = node558_l & pixel[93];
      node559_l = node558_l & ~pixel[93];
      node560 = node559_l;
      node561 = node559_r;
      node562_r = node558_r & pixel[329];
      node562_l = node558_r & ~pixel[329];
      node563 = node562_l;
      node564 = node562_r;
      node565_r = node557_r & pixel[268];
      node565_l = node557_r & ~pixel[268];
      node566_r = node565_l & pixel[230];
      node566_l = node565_l & ~pixel[230];
      node567 = node566_l;
      node568 = node566_r;
      node569_r = node565_r & pixel[248];
      node569_l = node565_r & ~pixel[248];
      node570 = node569_l;
      node571 = node569_r;
      node572_r = node556_r & pixel[304];
      node572_l = node556_r & ~pixel[304];
      node573_r = node572_l & pixel[464];
      node573_l = node572_l & ~pixel[464];
      node574_r = node573_l & pixel[574];
      node574_l = node573_l & ~pixel[574];
      node575 = node574_l;
      node576 = node574_r;
      node577_r = node573_r & pixel[267];
      node577_l = node573_r & ~pixel[267];
      node578 = node577_l;
      node579 = node577_r;
      node580_r = node572_r & pixel[295];
      node580_l = node572_r & ~pixel[295];
      node581 = node580_l;
      node582_r = node580_r & pixel[425];
      node582_l = node580_r & ~pixel[425];
      node583 = node582_l;
      node584 = node582_r;
      node585_r = node555_r & pixel[484];
      node585_l = node555_r & ~pixel[484];
      node586_r = node585_l & pixel[123];
      node586_l = node585_l & ~pixel[123];
      node587_r = node586_l & pixel[375];
      node587_l = node586_l & ~pixel[375];
      node588_r = node587_l & pixel[328];
      node588_l = node587_l & ~pixel[328];
      node589 = node588_l;
      node590 = node588_r;
      node591 = node587_r;
      node592 = node586_r;
      node593_r = node585_r & pixel[486];
      node593_l = node585_r & ~pixel[486];
      node594 = node593_l;
      node595_r = node593_r & pixel[436];
      node595_l = node593_r & ~pixel[436];
      node596 = node595_l;
      node597 = node595_r;
      node598_r = node554_r & pixel[270];
      node598_l = node554_r & ~pixel[270];
      node599_r = node598_l & pixel[354];
      node599_l = node598_l & ~pixel[354];
      node600_r = node599_l & pixel[188];
      node600_l = node599_l & ~pixel[188];
      node601_r = node600_l & pixel[236];
      node601_l = node600_l & ~pixel[236];
      node602_r = node601_l & pixel[208];
      node602_l = node601_l & ~pixel[208];
      node603 = node602_l;
      node604 = node602_r;
      node605_r = node601_r & pixel[455];
      node605_l = node601_r & ~pixel[455];
      node606 = node605_l;
      node607 = node605_r;
      node608_r = node600_r & pixel[275];
      node608_l = node600_r & ~pixel[275];
      node609_r = node608_l & pixel[300];
      node609_l = node608_l & ~pixel[300];
      node610 = node609_l;
      node611 = node609_r;
      node612_r = node608_r & pixel[385];
      node612_l = node608_r & ~pixel[385];
      node613 = node612_l;
      node614 = node612_r;
      node615_r = node599_r & pixel[526];
      node615_l = node599_r & ~pixel[526];
      node616_r = node615_l & pixel[192];
      node616_l = node615_l & ~pixel[192];
      node617_r = node616_l & pixel[436];
      node617_l = node616_l & ~pixel[436];
      node618 = node617_l;
      node619 = node617_r;
      node620_r = node616_r & pixel[187];
      node620_l = node616_r & ~pixel[187];
      node621 = node620_l;
      node622 = node620_r;
      node623_r = node615_r & pixel[285];
      node623_l = node615_r & ~pixel[285];
      node624_r = node623_l & pixel[545];
      node624_l = node623_l & ~pixel[545];
      node625 = node624_l;
      node626 = node624_r;
      node627_r = node623_r & pixel[201];
      node627_l = node623_r & ~pixel[201];
      node628 = node627_l;
      node629 = node627_r;
      node630_r = node598_r & pixel[383];
      node630_l = node598_r & ~pixel[383];
      node631_r = node630_l & pixel[681];
      node631_l = node630_l & ~pixel[681];
      node632_r = node631_l & pixel[298];
      node632_l = node631_l & ~pixel[298];
      node633_r = node632_l & pixel[655];
      node633_l = node632_l & ~pixel[655];
      node634 = node633_l;
      node635 = node633_r;
      node636_r = node632_r & pixel[154];
      node636_l = node632_r & ~pixel[154];
      node637 = node636_l;
      node638 = node636_r;
      node639_r = node631_r & pixel[659];
      node639_l = node631_r & ~pixel[659];
      node640_r = node639_l & pixel[549];
      node640_l = node639_l & ~pixel[549];
      node641 = node640_l;
      node642 = node640_r;
      node643_r = node639_r & pixel[454];
      node643_l = node639_r & ~pixel[454];
      node644 = node643_l;
      node645 = node643_r;
      node646_r = node630_r & pixel[155];
      node646_l = node630_r & ~pixel[155];
      node647_r = node646_l & pixel[431];
      node647_l = node646_l & ~pixel[431];
      node648_r = node647_l & pixel[245];
      node648_l = node647_l & ~pixel[245];
      node649 = node648_l;
      node650 = node648_r;
      node651_r = node647_r & pixel[498];
      node651_l = node647_r & ~pixel[498];
      node652 = node651_l;
      node653 = node651_r;
      node654_r = node646_r & pixel[235];
      node654_l = node646_r & ~pixel[235];
      node655_r = node654_l & pixel[567];
      node655_l = node654_l & ~pixel[567];
      node656 = node655_l;
      node657 = node655_r;
      node658_r = node654_r & pixel[553];
      node658_l = node654_r & ~pixel[553];
      node659 = node658_l;
      node660 = node658_r;
      node661_r = node427_r & pixel[685];
      node661_l = node427_r & ~pixel[685];
      node662_r = node661_l & pixel[217];
      node662_l = node661_l & ~pixel[217];
      node663_r = node662_l & pixel[214];
      node663_l = node662_l & ~pixel[214];
      node664_r = node663_l & pixel[663];
      node664_l = node663_l & ~pixel[663];
      node665_r = node664_l & pixel[296];
      node665_l = node664_l & ~pixel[296];
      node666_r = node665_l & pixel[241];
      node666_l = node665_l & ~pixel[241];
      node667_r = node666_l & pixel[661];
      node667_l = node666_l & ~pixel[661];
      node668 = node667_l;
      node669 = node667_r;
      node670_r = node666_r & pixel[659];
      node670_l = node666_r & ~pixel[659];
      node671 = node670_l;
      node672 = node670_r;
      node673_r = node665_r & pixel[414];
      node673_l = node665_r & ~pixel[414];
      node674_r = node673_l & pixel[375];
      node674_l = node673_l & ~pixel[375];
      node675 = node674_l;
      node676 = node674_r;
      node677_r = node673_r & pixel[485];
      node677_l = node673_r & ~pixel[485];
      node678 = node677_l;
      node679 = node677_r;
      node680_r = node664_r & pixel[373];
      node680_l = node664_r & ~pixel[373];
      node681_r = node680_l & pixel[404];
      node681_l = node680_l & ~pixel[404];
      node682_r = node681_l & pixel[608];
      node682_l = node681_l & ~pixel[608];
      node683 = node682_l;
      node684 = node682_r;
      node685_r = node681_r & pixel[497];
      node685_l = node681_r & ~pixel[497];
      node686 = node685_l;
      node687 = node685_r;
      node688_r = node680_r & pixel[602];
      node688_l = node680_r & ~pixel[602];
      node689_r = node688_l & pixel[384];
      node689_l = node688_l & ~pixel[384];
      node690 = node689_l;
      node691 = node689_r;
      node692_r = node688_r & pixel[342];
      node692_l = node688_r & ~pixel[342];
      node693 = node692_l;
      node694 = node692_r;
      node695_r = node663_r & pixel[461];
      node695_l = node663_r & ~pixel[461];
      node696_r = node695_l & pixel[378];
      node696_l = node695_l & ~pixel[378];
      node697_r = node696_l & pixel[180];
      node697_l = node696_l & ~pixel[180];
      node698_r = node697_l & pixel[271];
      node698_l = node697_l & ~pixel[271];
      node699 = node698_l;
      node700 = node698_r;
      node701_r = node697_r & pixel[601];
      node701_l = node697_r & ~pixel[601];
      node702 = node701_l;
      node703 = node701_r;
      node704_r = node696_r & pixel[180];
      node704_l = node696_r & ~pixel[180];
      node705_r = node704_l & pixel[293];
      node705_l = node704_l & ~pixel[293];
      node706 = node705_l;
      node707 = node705_r;
      node708_r = node704_r & pixel[464];
      node708_l = node704_r & ~pixel[464];
      node709 = node708_l;
      node710 = node708_r;
      node711_r = node695_r & pixel[298];
      node711_l = node695_r & ~pixel[298];
      node712_r = node711_l & pixel[574];
      node712_l = node711_l & ~pixel[574];
      node713_r = node712_l & pixel[454];
      node713_l = node712_l & ~pixel[454];
      node714 = node713_l;
      node715 = node713_r;
      node716_r = node712_r & pixel[549];
      node716_l = node712_r & ~pixel[549];
      node717 = node716_l;
      node718 = node716_r;
      node719_r = node711_r & pixel[601];
      node719_l = node711_r & ~pixel[601];
      node720_r = node719_l & pixel[183];
      node720_l = node719_l & ~pixel[183];
      node721 = node720_l;
      node722 = node720_r;
      node723_r = node719_r & pixel[546];
      node723_l = node719_r & ~pixel[546];
      node724 = node723_l;
      node725 = node723_r;
      node726_r = node662_r & pixel[213];
      node726_l = node662_r & ~pixel[213];
      node727_r = node726_l & pixel[158];
      node727_l = node726_l & ~pixel[158];
      node728_r = node727_l & pixel[296];
      node728_l = node727_l & ~pixel[296];
      node729_r = node728_l & pixel[488];
      node729_l = node728_l & ~pixel[488];
      node730 = node729_l;
      node731_r = node729_r & pixel[98];
      node731_l = node729_r & ~pixel[98];
      node732 = node731_l;
      node733 = node731_r;
      node734_r = node728_r & pixel[598];
      node734_l = node728_r & ~pixel[598];
      node735_r = node734_l & pixel[427];
      node735_l = node734_l & ~pixel[427];
      node736 = node735_l;
      node737 = node735_r;
      node738_r = node734_r & pixel[463];
      node738_l = node734_r & ~pixel[463];
      node739 = node738_l;
      node740 = node738_r;
      node741_r = node727_r & pixel[273];
      node741_l = node727_r & ~pixel[273];
      node742_r = node741_l & pixel[270];
      node742_l = node741_l & ~pixel[270];
      node743_r = node742_l & pixel[653];
      node743_l = node742_l & ~pixel[653];
      node744 = node743_l;
      node745 = node743_r;
      node746_r = node742_r & pixel[351];
      node746_l = node742_r & ~pixel[351];
      node747 = node746_l;
      node748 = node746_r;
      node749_r = node741_r & pixel[291];
      node749_l = node741_r & ~pixel[291];
      node750_r = node749_l & pixel[412];
      node750_l = node749_l & ~pixel[412];
      node751 = node750_l;
      node752 = node750_r;
      node753_r = node749_r & pixel[342];
      node753_l = node749_r & ~pixel[342];
      node754 = node753_l;
      node755 = node753_r;
      node756_r = node726_r & pixel[708];
      node756_l = node726_r & ~pixel[708];
      node757_r = node756_l & pixel[376];
      node757_l = node756_l & ~pixel[376];
      node758_r = node757_l & pixel[522];
      node758_l = node757_l & ~pixel[522];
      node759_r = node758_l & pixel[349];
      node759_l = node758_l & ~pixel[349];
      node760 = node759_l;
      node761 = node759_r;
      node762_r = node758_r & pixel[245];
      node762_l = node758_r & ~pixel[245];
      node763 = node762_l;
      node764 = node762_r;
      node765_r = node757_r & pixel[232];
      node765_l = node757_r & ~pixel[232];
      node766_r = node765_l & pixel[242];
      node766_l = node765_l & ~pixel[242];
      node767 = node766_l;
      node768 = node766_r;
      node769_r = node765_r & pixel[460];
      node769_l = node765_r & ~pixel[460];
      node770 = node769_l;
      node771 = node769_r;
      node772_r = node756_r & pixel[470];
      node772_l = node756_r & ~pixel[470];
      node773_r = node772_l & pixel[378];
      node773_l = node772_l & ~pixel[378];
      node774_r = node773_l & pixel[269];
      node774_l = node773_l & ~pixel[269];
      node775 = node774_l;
      node776 = node774_r;
      node777 = node773_r;
      node778 = node772_r;
      node779_r = node661_r & pixel[323];
      node779_l = node661_r & ~pixel[323];
      node780_r = node779_l & pixel[457];
      node780_l = node779_l & ~pixel[457];
      node781_r = node780_l & pixel[349];
      node781_l = node780_l & ~pixel[349];
      node782_r = node781_l & pixel[515];
      node782_l = node781_l & ~pixel[515];
      node783_r = node782_l & pixel[289];
      node783_l = node782_l & ~pixel[289];
      node784 = node783_l;
      node785_r = node783_r & pixel[467];
      node785_l = node783_r & ~pixel[467];
      node786 = node785_l;
      node787 = node785_r;
      node788_r = node782_r & pixel[468];
      node788_l = node782_r & ~pixel[468];
      node789_r = node788_l & pixel[609];
      node789_l = node788_l & ~pixel[609];
      node790 = node789_l;
      node791 = node789_r;
      node792_r = node788_r & pixel[463];
      node792_l = node788_r & ~pixel[463];
      node793 = node792_l;
      node794 = node792_r;
      node795_r = node781_r & pixel[515];
      node795_l = node781_r & ~pixel[515];
      node796 = node795_l;
      node797_r = node795_r & pixel[406];
      node797_l = node795_r & ~pixel[406];
      node798_r = node797_l & pixel[188];
      node798_l = node797_l & ~pixel[188];
      node799 = node798_l;
      node800 = node798_r;
      node801_r = node797_r & pixel[352];
      node801_l = node797_r & ~pixel[352];
      node802 = node801_l;
      node803 = node801_r;
      node804_r = node780_r & pixel[461];
      node804_l = node780_r & ~pixel[461];
      node805_r = node804_l & pixel[659];
      node805_l = node804_l & ~pixel[659];
      node806_r = node805_l & pixel[188];
      node806_l = node805_l & ~pixel[188];
      node807_r = node806_l & pixel[484];
      node807_l = node806_l & ~pixel[484];
      node808 = node807_l;
      node809 = node807_r;
      node810 = node806_r;
      node811_r = node805_r & pixel[515];
      node811_l = node805_r & ~pixel[515];
      node812_r = node811_l & pixel[186];
      node812_l = node811_l & ~pixel[186];
      node813 = node812_l;
      node814 = node812_r;
      node815_r = node811_r & pixel[629];
      node815_l = node811_r & ~pixel[629];
      node816 = node815_l;
      node817 = node815_r;
      node818_r = node804_r & pixel[404];
      node818_l = node804_r & ~pixel[404];
      node819_r = node818_l & pixel[243];
      node819_l = node818_l & ~pixel[243];
      node820_r = node819_l & pixel[183];
      node820_l = node819_l & ~pixel[183];
      node821 = node820_l;
      node822 = node820_r;
      node823_r = node819_r & pixel[437];
      node823_l = node819_r & ~pixel[437];
      node824 = node823_l;
      node825 = node823_r;
      node826_r = node818_r & pixel[598];
      node826_l = node818_r & ~pixel[598];
      node827_r = node826_l & pixel[375];
      node827_l = node826_l & ~pixel[375];
      node828 = node827_l;
      node829 = node827_r;
      node830_r = node826_r & pixel[376];
      node830_l = node826_r & ~pixel[376];
      node831 = node830_l;
      node832 = node830_r;
      node833_r = node779_r & pixel[455];
      node833_l = node779_r & ~pixel[455];
      node834_r = node833_l & pixel[384];
      node834_l = node833_l & ~pixel[384];
      node835_r = node834_l & pixel[217];
      node835_l = node834_l & ~pixel[217];
      node836_r = node835_l & pixel[468];
      node836_l = node835_l & ~pixel[468];
      node837_r = node836_l & pixel[406];
      node837_l = node836_l & ~pixel[406];
      node838 = node837_l;
      node839 = node837_r;
      node840_r = node836_r & pixel[493];
      node840_l = node836_r & ~pixel[493];
      node841 = node840_l;
      node842 = node840_r;
      node843_r = node835_r & pixel[431];
      node843_l = node835_r & ~pixel[431];
      node844 = node843_l;
      node845_r = node843_r & pixel[624];
      node845_l = node843_r & ~pixel[624];
      node846 = node845_l;
      node847 = node845_r;
      node848_r = node834_r & pixel[296];
      node848_l = node834_r & ~pixel[296];
      node849_r = node848_l & pixel[440];
      node849_l = node848_l & ~pixel[440];
      node850_r = node849_l & pixel[245];
      node850_l = node849_l & ~pixel[245];
      node851 = node850_l;
      node852 = node850_r;
      node853_r = node849_r & pixel[683];
      node853_l = node849_r & ~pixel[683];
      node854 = node853_l;
      node855 = node853_r;
      node856_r = node848_r & pixel[489];
      node856_l = node848_r & ~pixel[489];
      node857_r = node856_l & pixel[231];
      node857_l = node856_l & ~pixel[231];
      node858 = node857_l;
      node859 = node857_r;
      node860_r = node856_r & pixel[374];
      node860_l = node856_r & ~pixel[374];
      node861 = node860_l;
      node862 = node860_r;
      node863_r = node833_r & pixel[487];
      node863_l = node833_r & ~pixel[487];
      node864_r = node863_l & pixel[484];
      node864_l = node863_l & ~pixel[484];
      node865 = node864_l;
      node866 = node864_r;
      node867_r = node863_r & pixel[628];
      node867_l = node863_r & ~pixel[628];
      node868_r = node867_l & pixel[175];
      node868_l = node867_l & ~pixel[175];
      node869 = node868_l;
      node870_r = node868_r & pixel[190];
      node870_l = node868_r & ~pixel[190];
      node871 = node870_l;
      node872 = node870_r;
      node873_r = node867_r & pixel[635];
      node873_l = node867_r & ~pixel[635];
      node874_r = node873_l & pixel[471];
      node874_l = node873_l & ~pixel[471];
      node875 = node874_l;
      node876 = node874_r;
      node877_r = node873_r & pixel[379];
      node877_l = node873_r & ~pixel[379];
      node878 = node877_l;
      node879 = node877_r;
      node880_r = node0_r & pixel[359];
      node880_l = node0_r & ~pixel[359];
      node881_r = node880_l & pixel[412];
      node881_l = node880_l & ~pixel[412];
      node882_r = node881_l & pixel[376];
      node882_l = node881_l & ~pixel[376];
      node883_r = node882_l & pixel[551];
      node883_l = node882_l & ~pixel[551];
      node884_r = node883_l & pixel[436];
      node884_l = node883_l & ~pixel[436];
      node885_r = node884_l & pixel[405];
      node885_l = node884_l & ~pixel[405];
      node886_r = node885_l & pixel[487];
      node886_l = node885_l & ~pixel[487];
      node887_r = node886_l & pixel[653];
      node887_l = node886_l & ~pixel[653];
      node888_r = node887_l & pixel[460];
      node888_l = node887_l & ~pixel[460];
      node889 = node888_l;
      node890 = node888_r;
      node891_r = node887_r & pixel[323];
      node891_l = node887_r & ~pixel[323];
      node892 = node891_l;
      node893 = node891_r;
      node894_r = node886_r & pixel[152];
      node894_l = node886_r & ~pixel[152];
      node895_r = node894_l & pixel[408];
      node895_l = node894_l & ~pixel[408];
      node896 = node895_l;
      node897 = node895_r;
      node898_r = node894_r & pixel[345];
      node898_l = node894_r & ~pixel[345];
      node899 = node898_l;
      node900 = node898_r;
      node901_r = node885_r & pixel[180];
      node901_l = node885_r & ~pixel[180];
      node902_r = node901_l & pixel[629];
      node902_l = node901_l & ~pixel[629];
      node903_r = node902_l & pixel[293];
      node903_l = node902_l & ~pixel[293];
      node904 = node903_l;
      node905 = node903_r;
      node906_r = node902_r & pixel[124];
      node906_l = node902_r & ~pixel[124];
      node907 = node906_l;
      node908 = node906_r;
      node909_r = node901_r & pixel[293];
      node909_l = node901_r & ~pixel[293];
      node910_r = node909_l & pixel[548];
      node910_l = node909_l & ~pixel[548];
      node911 = node910_l;
      node912 = node910_r;
      node913_r = node909_r & pixel[498];
      node913_l = node909_r & ~pixel[498];
      node914 = node913_l;
      node915 = node913_r;
      node916_r = node884_r & pixel[605];
      node916_l = node884_r & ~pixel[605];
      node917_r = node916_l & pixel[152];
      node917_l = node916_l & ~pixel[152];
      node918_r = node917_l & pixel[706];
      node918_l = node917_l & ~pixel[706];
      node919_r = node918_l & pixel[574];
      node919_l = node918_l & ~pixel[574];
      node920 = node919_l;
      node921 = node919_r;
      node922_r = node918_r & pixel[598];
      node922_l = node918_r & ~pixel[598];
      node923 = node922_l;
      node924 = node922_r;
      node925_r = node917_r & pixel[321];
      node925_l = node917_r & ~pixel[321];
      node926_r = node925_l & pixel[346];
      node926_l = node925_l & ~pixel[346];
      node927 = node926_l;
      node928 = node926_r;
      node929_r = node925_r & pixel[328];
      node929_l = node925_r & ~pixel[328];
      node930 = node929_l;
      node931 = node929_r;
      node932_r = node916_r & pixel[655];
      node932_l = node916_r & ~pixel[655];
      node933_r = node932_l & pixel[467];
      node933_l = node932_l & ~pixel[467];
      node934_r = node933_l & pixel[373];
      node934_l = node933_l & ~pixel[373];
      node935 = node934_l;
      node936 = node934_r;
      node937_r = node933_r & pixel[580];
      node937_l = node933_r & ~pixel[580];
      node938 = node937_l;
      node939 = node937_r;
      node940_r = node932_r & pixel[550];
      node940_l = node932_r & ~pixel[550];
      node941_r = node940_l & pixel[549];
      node941_l = node940_l & ~pixel[549];
      node942 = node941_l;
      node943 = node941_r;
      node944_r = node940_r & pixel[327];
      node944_l = node940_r & ~pixel[327];
      node945 = node944_l;
      node946 = node944_r;
      node947_r = node883_r & pixel[659];
      node947_l = node883_r & ~pixel[659];
      node948_r = node947_l & pixel[461];
      node948_l = node947_l & ~pixel[461];
      node949_r = node948_l & pixel[515];
      node949_l = node948_l & ~pixel[515];
      node950_r = node949_l & pixel[629];
      node950_l = node949_l & ~pixel[629];
      node951_r = node950_l & pixel[541];
      node951_l = node950_l & ~pixel[541];
      node952 = node951_l;
      node953 = node951_r;
      node954_r = node950_r & pixel[353];
      node954_l = node950_r & ~pixel[353];
      node955 = node954_l;
      node956 = node954_r;
      node957_r = node949_r & pixel[293];
      node957_l = node949_r & ~pixel[293];
      node958_r = node957_l & pixel[236];
      node958_l = node957_l & ~pixel[236];
      node959 = node958_l;
      node960 = node958_r;
      node961_r = node957_r & pixel[235];
      node961_l = node957_r & ~pixel[235];
      node962 = node961_l;
      node963 = node961_r;
      node964_r = node948_r & pixel[390];
      node964_l = node948_r & ~pixel[390];
      node965_r = node964_l & pixel[400];
      node965_l = node964_l & ~pixel[400];
      node966_r = node965_l & pixel[346];
      node966_l = node965_l & ~pixel[346];
      node967 = node966_l;
      node968 = node966_r;
      node969_r = node965_r & pixel[520];
      node969_l = node965_r & ~pixel[520];
      node970 = node969_l;
      node971 = node969_r;
      node972 = node964_r;
      node973_r = node947_r & pixel[442];
      node973_l = node947_r & ~pixel[442];
      node974_r = node973_l & pixel[373];
      node974_l = node973_l & ~pixel[373];
      node975_r = node974_l & pixel[297];
      node975_l = node974_l & ~pixel[297];
      node976_r = node975_l & pixel[462];
      node976_l = node975_l & ~pixel[462];
      node977 = node976_l;
      node978 = node976_r;
      node979_r = node975_r & pixel[433];
      node979_l = node975_r & ~pixel[433];
      node980 = node979_l;
      node981 = node979_r;
      node982_r = node974_r & pixel[299];
      node982_l = node974_r & ~pixel[299];
      node983_r = node982_l & pixel[127];
      node983_l = node982_l & ~pixel[127];
      node984 = node983_l;
      node985 = node983_r;
      node986_r = node982_r & pixel[461];
      node986_l = node982_r & ~pixel[461];
      node987 = node986_l;
      node988 = node986_r;
      node989_r = node973_r & pixel[464];
      node989_l = node973_r & ~pixel[464];
      node990_r = node989_l & pixel[428];
      node990_l = node989_l & ~pixel[428];
      node991_r = node990_l & pixel[539];
      node991_l = node990_l & ~pixel[539];
      node992 = node991_l;
      node993 = node991_r;
      node994 = node990_r;
      node995 = node989_r;
      node996_r = node882_r & pixel[486];
      node996_l = node882_r & ~pixel[486];
      node997_r = node996_l & pixel[150];
      node997_l = node996_l & ~pixel[150];
      node998_r = node997_l & pixel[319];
      node998_l = node997_l & ~pixel[319];
      node999_r = node998_l & pixel[275];
      node999_l = node998_l & ~pixel[275];
      node1000_r = node999_l & pixel[455];
      node1000_l = node999_l & ~pixel[455];
      node1001_r = node1000_l & pixel[624];
      node1001_l = node1000_l & ~pixel[624];
      node1002 = node1001_l;
      node1003 = node1001_r;
      node1004_r = node1000_r & pixel[427];
      node1004_l = node1000_r & ~pixel[427];
      node1005 = node1004_l;
      node1006 = node1004_r;
      node1007_r = node999_r & pixel[384];
      node1007_l = node999_r & ~pixel[384];
      node1008_r = node1007_l & pixel[184];
      node1008_l = node1007_l & ~pixel[184];
      node1009 = node1008_l;
      node1010 = node1008_r;
      node1011_r = node1007_r & pixel[620];
      node1011_l = node1007_r & ~pixel[620];
      node1012 = node1011_l;
      node1013 = node1011_r;
      node1014_r = node998_r & pixel[328];
      node1014_l = node998_r & ~pixel[328];
      node1015_r = node1014_l & pixel[219];
      node1015_l = node1014_l & ~pixel[219];
      node1016_r = node1015_l & pixel[263];
      node1016_l = node1015_l & ~pixel[263];
      node1017 = node1016_l;
      node1018 = node1016_r;
      node1019_r = node1015_r & pixel[709];
      node1019_l = node1015_r & ~pixel[709];
      node1020 = node1019_l;
      node1021 = node1019_r;
      node1022_r = node1014_r & pixel[189];
      node1022_l = node1014_r & ~pixel[189];
      node1023_r = node1022_l & pixel[522];
      node1023_l = node1022_l & ~pixel[522];
      node1024 = node1023_l;
      node1025 = node1023_r;
      node1026_r = node1022_r & pixel[324];
      node1026_l = node1022_r & ~pixel[324];
      node1027 = node1026_l;
      node1028 = node1026_r;
      node1029_r = node997_r & pixel[316];
      node1029_l = node997_r & ~pixel[316];
      node1030_r = node1029_l & pixel[632];
      node1030_l = node1029_l & ~pixel[632];
      node1031_r = node1030_l & pixel[581];
      node1031_l = node1030_l & ~pixel[581];
      node1032_r = node1031_l & pixel[351];
      node1032_l = node1031_l & ~pixel[351];
      node1033 = node1032_l;
      node1034 = node1032_r;
      node1035_r = node1031_r & pixel[688];
      node1035_l = node1031_r & ~pixel[688];
      node1036 = node1035_l;
      node1037 = node1035_r;
      node1038_r = node1030_r & pixel[263];
      node1038_l = node1030_r & ~pixel[263];
      node1039_r = node1038_l & pixel[458];
      node1039_l = node1038_l & ~pixel[458];
      node1040 = node1039_l;
      node1041 = node1039_r;
      node1042_r = node1038_r & pixel[295];
      node1042_l = node1038_r & ~pixel[295];
      node1043 = node1042_l;
      node1044 = node1042_r;
      node1045_r = node1029_r & pixel[260];
      node1045_l = node1029_r & ~pixel[260];
      node1046_r = node1045_l & pixel[325];
      node1046_l = node1045_l & ~pixel[325];
      node1047_r = node1046_l & pixel[323];
      node1047_l = node1046_l & ~pixel[323];
      node1048 = node1047_l;
      node1049 = node1047_r;
      node1050_r = node1046_r & pixel[517];
      node1050_l = node1046_r & ~pixel[517];
      node1051 = node1050_l;
      node1052 = node1050_r;
      node1053_r = node1045_r & pixel[228];
      node1053_l = node1045_r & ~pixel[228];
      node1054_r = node1053_l & pixel[488];
      node1054_l = node1053_l & ~pixel[488];
      node1055 = node1054_l;
      node1056 = node1054_r;
      node1057_r = node1053_r & pixel[353];
      node1057_l = node1053_r & ~pixel[353];
      node1058 = node1057_l;
      node1059 = node1057_r;
      node1060_r = node996_r & pixel[299];
      node1060_l = node996_r & ~pixel[299];
      node1061_r = node1060_l & pixel[500];
      node1061_l = node1060_l & ~pixel[500];
      node1062_r = node1061_l & pixel[151];
      node1062_l = node1061_l & ~pixel[151];
      node1063_r = node1062_l & pixel[466];
      node1063_l = node1062_l & ~pixel[466];
      node1064_r = node1063_l & pixel[264];
      node1064_l = node1063_l & ~pixel[264];
      node1065 = node1064_l;
      node1066 = node1064_r;
      node1067_r = node1063_r & pixel[234];
      node1067_l = node1063_r & ~pixel[234];
      node1068 = node1067_l;
      node1069 = node1067_r;
      node1070_r = node1062_r & pixel[545];
      node1070_l = node1062_r & ~pixel[545];
      node1071_r = node1070_l & pixel[407];
      node1071_l = node1070_l & ~pixel[407];
      node1072 = node1071_l;
      node1073 = node1071_r;
      node1074_r = node1070_r & pixel[410];
      node1074_l = node1070_r & ~pixel[410];
      node1075 = node1074_l;
      node1076 = node1074_r;
      node1077_r = node1061_r & pixel[551];
      node1077_l = node1061_r & ~pixel[551];
      node1078_r = node1077_l & pixel[522];
      node1078_l = node1077_l & ~pixel[522];
      node1079_r = node1078_l & pixel[346];
      node1079_l = node1078_l & ~pixel[346];
      node1080 = node1079_l;
      node1081 = node1079_r;
      node1082_r = node1078_r & pixel[653];
      node1082_l = node1078_r & ~pixel[653];
      node1083 = node1082_l;
      node1084 = node1082_r;
      node1085_r = node1077_r & pixel[409];
      node1085_l = node1077_r & ~pixel[409];
      node1086 = node1085_l;
      node1087_r = node1085_r & pixel[178];
      node1087_l = node1085_r & ~pixel[178];
      node1088 = node1087_l;
      node1089 = node1087_r;
      node1090_r = node1060_r & pixel[554];
      node1090_l = node1060_r & ~pixel[554];
      node1091_r = node1090_l & pixel[210];
      node1091_l = node1090_l & ~pixel[210];
      node1092_r = node1091_l & pixel[207];
      node1092_l = node1091_l & ~pixel[207];
      node1093_r = node1092_l & pixel[292];
      node1093_l = node1092_l & ~pixel[292];
      node1094 = node1093_l;
      node1095 = node1093_r;
      node1096_r = node1092_r & pixel[638];
      node1096_l = node1092_r & ~pixel[638];
      node1097 = node1096_l;
      node1098 = node1096_r;
      node1099_r = node1091_r & pixel[380];
      node1099_l = node1091_r & ~pixel[380];
      node1100_r = node1099_l & pixel[438];
      node1100_l = node1099_l & ~pixel[438];
      node1101 = node1100_l;
      node1102 = node1100_r;
      node1103_r = node1099_r & pixel[508];
      node1103_l = node1099_r & ~pixel[508];
      node1104 = node1103_l;
      node1105 = node1103_r;
      node1106_r = node1090_r & pixel[371];
      node1106_l = node1090_r & ~pixel[371];
      node1107_r = node1106_l & pixel[483];
      node1107_l = node1106_l & ~pixel[483];
      node1108_r = node1107_l & pixel[318];
      node1108_l = node1107_l & ~pixel[318];
      node1109 = node1108_l;
      node1110 = node1108_r;
      node1111_r = node1107_r & pixel[660];
      node1111_l = node1107_r & ~pixel[660];
      node1112 = node1111_l;
      node1113 = node1111_r;
      node1114_r = node1106_r & pixel[426];
      node1114_l = node1106_r & ~pixel[426];
      node1115 = node1114_l;
      node1116_r = node1114_r & pixel[128];
      node1116_l = node1114_r & ~pixel[128];
      node1117 = node1116_l;
      node1118 = node1116_r;
      node1119_r = node881_r & pixel[462];
      node1119_l = node881_r & ~pixel[462];
      node1120_r = node1119_l & pixel[350];
      node1120_l = node1119_l & ~pixel[350];
      node1121_r = node1120_l & pixel[372];
      node1121_l = node1120_l & ~pixel[372];
      node1122_r = node1121_l & pixel[516];
      node1122_l = node1121_l & ~pixel[516];
      node1123_r = node1122_l & pixel[352];
      node1123_l = node1122_l & ~pixel[352];
      node1124_r = node1123_l & pixel[379];
      node1124_l = node1123_l & ~pixel[379];
      node1125_r = node1124_l & pixel[457];
      node1125_l = node1124_l & ~pixel[457];
      node1126 = node1125_l;
      node1127 = node1125_r;
      node1128_r = node1124_r & pixel[521];
      node1128_l = node1124_r & ~pixel[521];
      node1129 = node1128_l;
      node1130 = node1128_r;
      node1131_r = node1123_r & pixel[151];
      node1131_l = node1123_r & ~pixel[151];
      node1132_r = node1131_l & pixel[431];
      node1132_l = node1131_l & ~pixel[431];
      node1133 = node1132_l;
      node1134 = node1132_r;
      node1135_r = node1131_r & pixel[383];
      node1135_l = node1131_r & ~pixel[383];
      node1136 = node1135_l;
      node1137 = node1135_r;
      node1138_r = node1122_r & pixel[376];
      node1138_l = node1122_r & ~pixel[376];
      node1139_r = node1138_l & pixel[395];
      node1139_l = node1138_l & ~pixel[395];
      node1140_r = node1139_l & pixel[348];
      node1140_l = node1139_l & ~pixel[348];
      node1141 = node1140_l;
      node1142 = node1140_r;
      node1143_r = node1139_r & pixel[286];
      node1143_l = node1139_r & ~pixel[286];
      node1144 = node1143_l;
      node1145 = node1143_r;
      node1146_r = node1138_r & pixel[293];
      node1146_l = node1138_r & ~pixel[293];
      node1147 = node1146_l;
      node1148_r = node1146_r & pixel[177];
      node1148_l = node1146_r & ~pixel[177];
      node1149 = node1148_l;
      node1150 = node1148_r;
      node1151_r = node1121_r & pixel[405];
      node1151_l = node1121_r & ~pixel[405];
      node1152_r = node1151_l & pixel[185];
      node1152_l = node1151_l & ~pixel[185];
      node1153_r = node1152_l & pixel[240];
      node1153_l = node1152_l & ~pixel[240];
      node1154_r = node1153_l & pixel[596];
      node1154_l = node1153_l & ~pixel[596];
      node1155 = node1154_l;
      node1156 = node1154_r;
      node1157_r = node1153_r & pixel[384];
      node1157_l = node1153_r & ~pixel[384];
      node1158 = node1157_l;
      node1159 = node1157_r;
      node1160_r = node1152_r & pixel[73];
      node1160_l = node1152_r & ~pixel[73];
      node1161_r = node1160_l & pixel[99];
      node1161_l = node1160_l & ~pixel[99];
      node1162 = node1161_l;
      node1163 = node1161_r;
      node1164 = node1160_r;
      node1165_r = node1151_r & pixel[514];
      node1165_l = node1151_r & ~pixel[514];
      node1166_r = node1165_l & pixel[463];
      node1166_l = node1165_l & ~pixel[463];
      node1167_r = node1166_l & pixel[460];
      node1167_l = node1166_l & ~pixel[460];
      node1168 = node1167_l;
      node1169 = node1167_r;
      node1170_r = node1166_r & pixel[688];
      node1170_l = node1166_r & ~pixel[688];
      node1171 = node1170_l;
      node1172 = node1170_r;
      node1173_r = node1165_r & pixel[242];
      node1173_l = node1165_r & ~pixel[242];
      node1174 = node1173_l;
      node1175_r = node1173_r & pixel[327];
      node1175_l = node1173_r & ~pixel[327];
      node1176 = node1175_l;
      node1177 = node1175_r;
      node1178_r = node1120_r & pixel[269];
      node1178_l = node1120_r & ~pixel[269];
      node1179_r = node1178_l & pixel[428];
      node1179_l = node1178_l & ~pixel[428];
      node1180_r = node1179_l & pixel[261];
      node1180_l = node1179_l & ~pixel[261];
      node1181_r = node1180_l & pixel[130];
      node1181_l = node1180_l & ~pixel[130];
      node1182_r = node1181_l & pixel[291];
      node1182_l = node1181_l & ~pixel[291];
      node1183 = node1182_l;
      node1184 = node1182_r;
      node1185_r = node1181_r & pixel[458];
      node1185_l = node1181_r & ~pixel[458];
      node1186 = node1185_l;
      node1187 = node1185_r;
      node1188_r = node1180_r & pixel[288];
      node1188_l = node1180_r & ~pixel[288];
      node1189_r = node1188_l & pixel[271];
      node1189_l = node1188_l & ~pixel[271];
      node1190 = node1189_l;
      node1191 = node1189_r;
      node1192_r = node1188_r & pixel[556];
      node1192_l = node1188_r & ~pixel[556];
      node1193 = node1192_l;
      node1194 = node1192_r;
      node1195_r = node1179_r & pixel[655];
      node1195_l = node1179_r & ~pixel[655];
      node1196_r = node1195_l & pixel[244];
      node1196_l = node1195_l & ~pixel[244];
      node1197_r = node1196_l & pixel[541];
      node1197_l = node1196_l & ~pixel[541];
      node1198 = node1197_l;
      node1199 = node1197_r;
      node1200_r = node1196_r & pixel[604];
      node1200_l = node1196_r & ~pixel[604];
      node1201 = node1200_l;
      node1202 = node1200_r;
      node1203_r = node1195_r & pixel[302];
      node1203_l = node1195_r & ~pixel[302];
      node1204_r = node1203_l & pixel[272];
      node1204_l = node1203_l & ~pixel[272];
      node1205 = node1204_l;
      node1206 = node1204_r;
      node1207_r = node1203_r & pixel[378];
      node1207_l = node1203_r & ~pixel[378];
      node1208 = node1207_l;
      node1209 = node1207_r;
      node1210_r = node1178_r & pixel[273];
      node1210_l = node1178_r & ~pixel[273];
      node1211_r = node1210_l & pixel[289];
      node1211_l = node1210_l & ~pixel[289];
      node1212_r = node1211_l & pixel[429];
      node1212_l = node1211_l & ~pixel[429];
      node1213_r = node1212_l & pixel[193];
      node1213_l = node1212_l & ~pixel[193];
      node1214 = node1213_l;
      node1215 = node1213_r;
      node1216_r = node1212_r & pixel[578];
      node1216_l = node1212_r & ~pixel[578];
      node1217 = node1216_l;
      node1218 = node1216_r;
      node1219_r = node1211_r & pixel[373];
      node1219_l = node1211_r & ~pixel[373];
      node1220_r = node1219_l & pixel[183];
      node1220_l = node1219_l & ~pixel[183];
      node1221 = node1220_l;
      node1222 = node1220_r;
      node1223_r = node1219_r & pixel[456];
      node1223_l = node1219_r & ~pixel[456];
      node1224 = node1223_l;
      node1225 = node1223_r;
      node1226_r = node1210_r & pixel[385];
      node1226_l = node1210_r & ~pixel[385];
      node1227_r = node1226_l & pixel[378];
      node1227_l = node1226_l & ~pixel[378];
      node1228_r = node1227_l & pixel[625];
      node1228_l = node1227_l & ~pixel[625];
      node1229 = node1228_l;
      node1230 = node1228_r;
      node1231_r = node1227_r & pixel[323];
      node1231_l = node1227_r & ~pixel[323];
      node1232 = node1231_l;
      node1233 = node1231_r;
      node1234_r = node1226_r & pixel[330];
      node1234_l = node1226_r & ~pixel[330];
      node1235_r = node1234_l & pixel[353];
      node1235_l = node1234_l & ~pixel[353];
      node1236 = node1235_l;
      node1237 = node1235_r;
      node1238_r = node1234_r & pixel[341];
      node1238_l = node1234_r & ~pixel[341];
      node1239 = node1238_l;
      node1240 = node1238_r;
      node1241_r = node1119_r & pixel[272];
      node1241_l = node1119_r & ~pixel[272];
      node1242_r = node1241_l & pixel[269];
      node1242_l = node1241_l & ~pixel[269];
      node1243_r = node1242_l & pixel[611];
      node1243_l = node1242_l & ~pixel[611];
      node1244_r = node1243_l & pixel[573];
      node1244_l = node1243_l & ~pixel[573];
      node1245_r = node1244_l & pixel[629];
      node1245_l = node1244_l & ~pixel[629];
      node1246_r = node1245_l & pixel[345];
      node1246_l = node1245_l & ~pixel[345];
      node1247 = node1246_l;
      node1248 = node1246_r;
      node1249_r = node1245_r & pixel[357];
      node1249_l = node1245_r & ~pixel[357];
      node1250 = node1249_l;
      node1251 = node1249_r;
      node1252_r = node1244_r & pixel[189];
      node1252_l = node1244_r & ~pixel[189];
      node1253_r = node1252_l & pixel[445];
      node1253_l = node1252_l & ~pixel[445];
      node1254 = node1253_l;
      node1255 = node1253_r;
      node1256_r = node1252_r & pixel[627];
      node1256_l = node1252_r & ~pixel[627];
      node1257 = node1256_l;
      node1258 = node1256_r;
      node1259_r = node1243_r & pixel[659];
      node1259_l = node1243_r & ~pixel[659];
      node1260_r = node1259_l & pixel[354];
      node1260_l = node1259_l & ~pixel[354];
      node1261 = node1260_l;
      node1262_r = node1260_r & pixel[669];
      node1262_l = node1260_r & ~pixel[669];
      node1263 = node1262_l;
      node1264 = node1262_r;
      node1265 = node1259_r;
      node1266_r = node1242_r & pixel[161];
      node1266_l = node1242_r & ~pixel[161];
      node1267_r = node1266_l & pixel[350];
      node1267_l = node1266_l & ~pixel[350];
      node1268_r = node1267_l & pixel[347];
      node1268_l = node1267_l & ~pixel[347];
      node1269_r = node1268_l & pixel[371];
      node1269_l = node1268_l & ~pixel[371];
      node1270 = node1269_l;
      node1271 = node1269_r;
      node1272_r = node1268_r & pixel[156];
      node1272_l = node1268_r & ~pixel[156];
      node1273 = node1272_l;
      node1274 = node1272_r;
      node1275_r = node1267_r & pixel[103];
      node1275_l = node1267_r & ~pixel[103];
      node1276_r = node1275_l & pixel[628];
      node1276_l = node1275_l & ~pixel[628];
      node1277 = node1276_l;
      node1278 = node1276_r;
      node1279 = node1275_r;
      node1280_r = node1266_r & pixel[294];
      node1280_l = node1266_r & ~pixel[294];
      node1281_r = node1280_l & pixel[565];
      node1281_l = node1280_l & ~pixel[565];
      node1282 = node1281_l;
      node1283_r = node1281_r & pixel[631];
      node1283_l = node1281_r & ~pixel[631];
      node1284 = node1283_l;
      node1285 = node1283_r;
      node1286_r = node1280_r & pixel[302];
      node1286_l = node1280_r & ~pixel[302];
      node1287_r = node1286_l & pixel[522];
      node1287_l = node1286_l & ~pixel[522];
      node1288 = node1287_l;
      node1289 = node1287_r;
      node1290_r = node1286_r & pixel[371];
      node1290_l = node1286_r & ~pixel[371];
      node1291 = node1290_l;
      node1292 = node1290_r;
      node1293_r = node1241_r & pixel[320];
      node1293_l = node1241_r & ~pixel[320];
      node1294_r = node1293_l & pixel[686];
      node1294_l = node1293_l & ~pixel[686];
      node1295_r = node1294_l & pixel[158];
      node1295_l = node1294_l & ~pixel[158];
      node1296_r = node1295_l & pixel[380];
      node1296_l = node1295_l & ~pixel[380];
      node1297_r = node1296_l & pixel[316];
      node1297_l = node1296_l & ~pixel[316];
      node1298 = node1297_l;
      node1299 = node1297_r;
      node1300_r = node1296_r & pixel[317];
      node1300_l = node1296_r & ~pixel[317];
      node1301 = node1300_l;
      node1302 = node1300_r;
      node1303_r = node1295_r & pixel[349];
      node1303_l = node1295_r & ~pixel[349];
      node1304_r = node1303_l & pixel[317];
      node1304_l = node1303_l & ~pixel[317];
      node1305 = node1304_l;
      node1306 = node1304_r;
      node1307_r = node1303_r & pixel[454];
      node1307_l = node1303_r & ~pixel[454];
      node1308 = node1307_l;
      node1309 = node1307_r;
      node1310_r = node1294_r & pixel[461];
      node1310_l = node1294_r & ~pixel[461];
      node1311_r = node1310_l & pixel[596];
      node1311_l = node1310_l & ~pixel[596];
      node1312 = node1311_l;
      node1313_r = node1311_r & pixel[552];
      node1313_l = node1311_r & ~pixel[552];
      node1314 = node1313_l;
      node1315 = node1313_r;
      node1316_r = node1310_r & pixel[316];
      node1316_l = node1310_r & ~pixel[316];
      node1317_r = node1316_l & pixel[581];
      node1317_l = node1316_l & ~pixel[581];
      node1318 = node1317_l;
      node1319 = node1317_r;
      node1320_r = node1316_r & pixel[415];
      node1320_l = node1316_r & ~pixel[415];
      node1321 = node1320_l;
      node1322 = node1320_r;
      node1323_r = node1293_r & pixel[406];
      node1323_l = node1293_r & ~pixel[406];
      node1324_r = node1323_l & pixel[453];
      node1324_l = node1323_l & ~pixel[453];
      node1325_r = node1324_l & pixel[400];
      node1325_l = node1324_l & ~pixel[400];
      node1326_r = node1325_l & pixel[374];
      node1326_l = node1325_l & ~pixel[374];
      node1327 = node1326_l;
      node1328 = node1326_r;
      node1329_r = node1325_r & pixel[484];
      node1329_l = node1325_r & ~pixel[484];
      node1330 = node1329_l;
      node1331 = node1329_r;
      node1332_r = node1324_r & pixel[715];
      node1332_l = node1324_r & ~pixel[715];
      node1333 = node1332_l;
      node1334 = node1332_r;
      node1335_r = node1323_r & pixel[655];
      node1335_l = node1323_r & ~pixel[655];
      node1336_r = node1335_l & pixel[522];
      node1336_l = node1335_l & ~pixel[522];
      node1337_r = node1336_l & pixel[213];
      node1337_l = node1336_l & ~pixel[213];
      node1338 = node1337_l;
      node1339 = node1337_r;
      node1340_r = node1336_r & pixel[453];
      node1340_l = node1336_r & ~pixel[453];
      node1341 = node1340_l;
      node1342 = node1340_r;
      node1343_r = node1335_r & pixel[707];
      node1343_l = node1335_r & ~pixel[707];
      node1344_r = node1343_l & pixel[515];
      node1344_l = node1343_l & ~pixel[515];
      node1345 = node1344_l;
      node1346 = node1344_r;
      node1347_r = node1343_r & pixel[248];
      node1347_l = node1343_r & ~pixel[248];
      node1348 = node1347_l;
      node1349 = node1347_r;
      node1350_r = node880_r & pixel[408];
      node1350_l = node880_r & ~pixel[408];
      node1351_r = node1350_l & pixel[399];
      node1351_l = node1350_l & ~pixel[399];
      node1352_r = node1351_l & pixel[151];
      node1352_l = node1351_l & ~pixel[151];
      node1353_r = node1352_l & pixel[492];
      node1353_l = node1352_l & ~pixel[492];
      node1354_r = node1353_l & pixel[333];
      node1354_l = node1353_l & ~pixel[333];
      node1355_r = node1354_l & pixel[414];
      node1355_l = node1354_l & ~pixel[414];
      node1356_r = node1355_l & pixel[290];
      node1356_l = node1355_l & ~pixel[290];
      node1357_r = node1356_l & pixel[579];
      node1357_l = node1356_l & ~pixel[579];
      node1358 = node1357_l;
      node1359 = node1357_r;
      node1360_r = node1356_r & pixel[511];
      node1360_l = node1356_r & ~pixel[511];
      node1361 = node1360_l;
      node1362 = node1360_r;
      node1363_r = node1355_r & pixel[214];
      node1363_l = node1355_r & ~pixel[214];
      node1364_r = node1363_l & pixel[378];
      node1364_l = node1363_l & ~pixel[378];
      node1365 = node1364_l;
      node1366 = node1364_r;
      node1367 = node1363_r;
      node1368 = node1354_r;
      node1369_r = node1353_r & pixel[188];
      node1369_l = node1353_r & ~pixel[188];
      node1370_r = node1369_l & pixel[322];
      node1370_l = node1369_l & ~pixel[322];
      node1371_r = node1370_l & pixel[318];
      node1371_l = node1370_l & ~pixel[318];
      node1372_r = node1371_l & pixel[378];
      node1372_l = node1371_l & ~pixel[378];
      node1373 = node1372_l;
      node1374 = node1372_r;
      node1375 = node1371_r;
      node1376_r = node1370_r & pixel[463];
      node1376_l = node1370_r & ~pixel[463];
      node1377 = node1376_l;
      node1378_r = node1376_r & pixel[385];
      node1378_l = node1376_r & ~pixel[385];
      node1379 = node1378_l;
      node1380 = node1378_r;
      node1381_r = node1369_r & pixel[607];
      node1381_l = node1369_r & ~pixel[607];
      node1382_r = node1381_l & pixel[553];
      node1382_l = node1381_l & ~pixel[553];
      node1383_r = node1382_l & pixel[483];
      node1383_l = node1382_l & ~pixel[483];
      node1384 = node1383_l;
      node1385 = node1383_r;
      node1386_r = node1382_r & pixel[269];
      node1386_l = node1382_r & ~pixel[269];
      node1387 = node1386_l;
      node1388 = node1386_r;
      node1389 = node1381_r;
      node1390_r = node1352_r & pixel[520];
      node1390_l = node1352_r & ~pixel[520];
      node1391_r = node1390_l & pixel[383];
      node1391_l = node1390_l & ~pixel[383];
      node1392_r = node1391_l & pixel[436];
      node1392_l = node1391_l & ~pixel[436];
      node1393_r = node1392_l & pixel[213];
      node1393_l = node1392_l & ~pixel[213];
      node1394_r = node1393_l & pixel[544];
      node1394_l = node1393_l & ~pixel[544];
      node1395 = node1394_l;
      node1396 = node1394_r;
      node1397 = node1393_r;
      node1398 = node1392_r;
      node1399_r = node1391_r & pixel[634];
      node1399_l = node1391_r & ~pixel[634];
      node1400 = node1399_l;
      node1401 = node1399_r;
      node1402_r = node1390_r & pixel[470];
      node1402_l = node1390_r & ~pixel[470];
      node1403_r = node1402_l & pixel[658];
      node1403_l = node1402_l & ~pixel[658];
      node1404 = node1403_l;
      node1405_r = node1403_r & pixel[360];
      node1405_l = node1403_r & ~pixel[360];
      node1406_r = node1405_l & pixel[328];
      node1406_l = node1405_l & ~pixel[328];
      node1407 = node1406_l;
      node1408 = node1406_r;
      node1409 = node1405_r;
      node1410_r = node1402_r & pixel[266];
      node1410_l = node1402_r & ~pixel[266];
      node1411_r = node1410_l & pixel[172];
      node1411_l = node1410_l & ~pixel[172];
      node1412 = node1411_l;
      node1413_r = node1411_r & pixel[213];
      node1413_l = node1411_r & ~pixel[213];
      node1414 = node1413_l;
      node1415 = node1413_r;
      node1416_r = node1410_r & pixel[370];
      node1416_l = node1410_r & ~pixel[370];
      node1417_r = node1416_l & pixel[543];
      node1417_l = node1416_l & ~pixel[543];
      node1418 = node1417_l;
      node1419 = node1417_r;
      node1420 = node1416_r;
      node1421_r = node1351_r & pixel[67];
      node1421_l = node1351_r & ~pixel[67];
      node1422_r = node1421_l & pixel[210];
      node1422_l = node1421_l & ~pixel[210];
      node1423_r = node1422_l & pixel[378];
      node1423_l = node1422_l & ~pixel[378];
      node1424_r = node1423_l & pixel[93];
      node1424_l = node1423_l & ~pixel[93];
      node1425_r = node1424_l & pixel[463];
      node1425_l = node1424_l & ~pixel[463];
      node1426_r = node1425_l & pixel[437];
      node1426_l = node1425_l & ~pixel[437];
      node1427 = node1426_l;
      node1428 = node1426_r;
      node1429_r = node1425_r & pixel[481];
      node1429_l = node1425_r & ~pixel[481];
      node1430 = node1429_l;
      node1431 = node1429_r;
      node1432_r = node1424_r & pixel[174];
      node1432_l = node1424_r & ~pixel[174];
      node1433_r = node1432_l & pixel[126];
      node1433_l = node1432_l & ~pixel[126];
      node1434 = node1433_l;
      node1435 = node1433_r;
      node1436 = node1432_r;
      node1437_r = node1423_r & pixel[215];
      node1437_l = node1423_r & ~pixel[215];
      node1438_r = node1437_l & pixel[415];
      node1438_l = node1437_l & ~pixel[415];
      node1439 = node1438_l;
      node1440_r = node1438_r & pixel[410];
      node1440_l = node1438_r & ~pixel[410];
      node1441 = node1440_l;
      node1442 = node1440_r;
      node1443_r = node1437_r & pixel[259];
      node1443_l = node1437_r & ~pixel[259];
      node1444 = node1443_l;
      node1445_r = node1443_r & pixel[578];
      node1445_l = node1443_r & ~pixel[578];
      node1446 = node1445_l;
      node1447 = node1445_r;
      node1448_r = node1422_r & pixel[244];
      node1448_l = node1422_r & ~pixel[244];
      node1449_r = node1448_l & pixel[350];
      node1449_l = node1448_l & ~pixel[350];
      node1450_r = node1449_l & pixel[188];
      node1450_l = node1449_l & ~pixel[188];
      node1451_r = node1450_l & pixel[329];
      node1451_l = node1450_l & ~pixel[329];
      node1452 = node1451_l;
      node1453 = node1451_r;
      node1454 = node1450_r;
      node1455_r = node1449_r & pixel[230];
      node1455_l = node1449_r & ~pixel[230];
      node1456_r = node1455_l & pixel[240];
      node1456_l = node1455_l & ~pixel[240];
      node1457 = node1456_l;
      node1458 = node1456_r;
      node1459 = node1455_r;
      node1460_r = node1448_r & pixel[405];
      node1460_l = node1448_r & ~pixel[405];
      node1461_r = node1460_l & pixel[273];
      node1461_l = node1460_l & ~pixel[273];
      node1462_r = node1461_l & pixel[313];
      node1462_l = node1461_l & ~pixel[313];
      node1463 = node1462_l;
      node1464 = node1462_r;
      node1465_r = node1461_r & pixel[344];
      node1465_l = node1461_r & ~pixel[344];
      node1466 = node1465_l;
      node1467 = node1465_r;
      node1468_r = node1460_r & pixel[344];
      node1468_l = node1460_r & ~pixel[344];
      node1469_r = node1468_l & pixel[182];
      node1469_l = node1468_l & ~pixel[182];
      node1470 = node1469_l;
      node1471 = node1469_r;
      node1472_r = node1468_r & pixel[501];
      node1472_l = node1468_r & ~pixel[501];
      node1473 = node1472_l;
      node1474 = node1472_r;
      node1475 = node1421_r;
      node1476_r = node1350_r & pixel[414];
      node1476_l = node1350_r & ~pixel[414];
      node1477_r = node1476_l & pixel[459];
      node1477_l = node1476_l & ~pixel[459];
      node1478_r = node1477_l & pixel[626];
      node1478_l = node1477_l & ~pixel[626];
      node1479_r = node1478_l & pixel[376];
      node1479_l = node1478_l & ~pixel[376];
      node1480_r = node1479_l & pixel[390];
      node1480_l = node1479_l & ~pixel[390];
      node1481 = node1480_l;
      node1482 = node1480_r;
      node1483_r = node1479_r & pixel[518];
      node1483_l = node1479_r & ~pixel[518];
      node1484 = node1483_l;
      node1485 = node1483_r;
      node1486_r = node1478_r & pixel[404];
      node1486_l = node1478_r & ~pixel[404];
      node1487_r = node1486_l & pixel[378];
      node1487_l = node1486_l & ~pixel[378];
      node1488_r = node1487_l & pixel[429];
      node1488_l = node1487_l & ~pixel[429];
      node1489 = node1488_l;
      node1490 = node1488_r;
      node1491_r = node1487_r & pixel[410];
      node1491_l = node1487_r & ~pixel[410];
      node1492 = node1491_l;
      node1493 = node1491_r;
      node1494_r = node1486_r & pixel[524];
      node1494_l = node1486_r & ~pixel[524];
      node1495_r = node1494_l & pixel[412];
      node1495_l = node1494_l & ~pixel[412];
      node1496_r = node1495_l & pixel[352];
      node1496_l = node1495_l & ~pixel[352];
      node1497 = node1496_l;
      node1498 = node1496_r;
      node1499_r = node1495_r & pixel[600];
      node1499_l = node1495_r & ~pixel[600];
      node1500 = node1499_l;
      node1501 = node1499_r;
      node1502_r = node1494_r & pixel[342];
      node1502_l = node1494_r & ~pixel[342];
      node1503 = node1502_l;
      node1504_r = node1502_r & pixel[580];
      node1504_l = node1502_r & ~pixel[580];
      node1505 = node1504_l;
      node1506 = node1504_r;
      node1507_r = node1477_r & pixel[466];
      node1507_l = node1477_r & ~pixel[466];
      node1508_r = node1507_l & pixel[735];
      node1508_l = node1507_l & ~pixel[735];
      node1509_r = node1508_l & pixel[215];
      node1509_l = node1508_l & ~pixel[215];
      node1510_r = node1509_l & pixel[398];
      node1510_l = node1509_l & ~pixel[398];
      node1511_r = node1510_l & pixel[209];
      node1511_l = node1510_l & ~pixel[209];
      node1512 = node1511_l;
      node1513 = node1511_r;
      node1514 = node1510_r;
      node1515 = node1509_r;
      node1516_r = node1508_r & pixel[706];
      node1516_l = node1508_r & ~pixel[706];
      node1517 = node1516_l;
      node1518 = node1516_r;
      node1519_r = node1507_r & pixel[482];
      node1519_l = node1507_r & ~pixel[482];
      node1520_r = node1519_l & pixel[572];
      node1520_l = node1519_l & ~pixel[572];
      node1521 = node1520_l;
      node1522_r = node1520_r & pixel[517];
      node1522_l = node1520_r & ~pixel[517];
      node1523 = node1522_l;
      node1524_r = node1522_r & pixel[286];
      node1524_l = node1522_r & ~pixel[286];
      node1525 = node1524_l;
      node1526 = node1524_r;
      node1527_r = node1519_r & pixel[242];
      node1527_l = node1519_r & ~pixel[242];
      node1528 = node1527_l;
      node1529_r = node1527_r & pixel[323];
      node1529_l = node1527_r & ~pixel[323];
      node1530 = node1529_l;
      node1531 = node1529_r;
      node1532_r = node1476_r & pixel[496];
      node1532_l = node1476_r & ~pixel[496];
      node1533_r = node1532_l & pixel[375];
      node1533_l = node1532_l & ~pixel[375];
      node1534_r = node1533_l & pixel[260];
      node1534_l = node1533_l & ~pixel[260];
      node1535_r = node1534_l & pixel[626];
      node1535_l = node1534_l & ~pixel[626];
      node1536_r = node1535_l & pixel[432];
      node1536_l = node1535_l & ~pixel[432];
      node1537_r = node1536_l & pixel[269];
      node1537_l = node1536_l & ~pixel[269];
      node1538 = node1537_l;
      node1539 = node1537_r;
      node1540_r = node1536_r & pixel[242];
      node1540_l = node1536_r & ~pixel[242];
      node1541 = node1540_l;
      node1542 = node1540_r;
      node1543 = node1535_r;
      node1544_r = node1534_r & pixel[695];
      node1544_l = node1534_r & ~pixel[695];
      node1545_r = node1544_l & pixel[579];
      node1545_l = node1544_l & ~pixel[579];
      node1546_r = node1545_l & pixel[178];
      node1546_l = node1545_l & ~pixel[178];
      node1547 = node1546_l;
      node1548 = node1546_r;
      node1549 = node1545_r;
      node1550 = node1544_r;
      node1551_r = node1533_r & pixel[443];
      node1551_l = node1533_r & ~pixel[443];
      node1552_r = node1551_l & pixel[129];
      node1552_l = node1551_l & ~pixel[129];
      node1553_r = node1552_l & pixel[655];
      node1553_l = node1552_l & ~pixel[655];
      node1554_r = node1553_l & pixel[567];
      node1554_l = node1553_l & ~pixel[567];
      node1555 = node1554_l;
      node1556 = node1554_r;
      node1557 = node1553_r;
      node1558_r = node1552_r & pixel[179];
      node1558_l = node1552_r & ~pixel[179];
      node1559 = node1558_l;
      node1560 = node1558_r;
      node1561_r = node1551_r & pixel[598];
      node1561_l = node1551_r & ~pixel[598];
      node1562_r = node1561_l & pixel[343];
      node1562_l = node1561_l & ~pixel[343];
      node1563 = node1562_l;
      node1564 = node1562_r;
      node1565_r = node1561_r & pixel[217];
      node1565_l = node1561_r & ~pixel[217];
      node1566_r = node1565_l & pixel[352];
      node1566_l = node1565_l & ~pixel[352];
      node1567 = node1566_l;
      node1568 = node1566_r;
      node1569 = node1565_r;
      node1570_r = node1532_r & pixel[240];
      node1570_l = node1532_r & ~pixel[240];
      node1571_r = node1570_l & pixel[189];
      node1571_l = node1570_l & ~pixel[189];
      node1572_r = node1571_l & pixel[653];
      node1572_l = node1571_l & ~pixel[653];
      node1573_r = node1572_l & pixel[635];
      node1573_l = node1572_l & ~pixel[635];
      node1574_r = node1573_l & pixel[576];
      node1574_l = node1573_l & ~pixel[576];
      node1575 = node1574_l;
      node1576 = node1574_r;
      node1577_r = node1573_r & pixel[443];
      node1577_l = node1573_r & ~pixel[443];
      node1578 = node1577_l;
      node1579 = node1577_r;
      node1580_r = node1572_r & pixel[378];
      node1580_l = node1572_r & ~pixel[378];
      node1581_r = node1580_l & pixel[230];
      node1581_l = node1580_l & ~pixel[230];
      node1582 = node1581_l;
      node1583 = node1581_r;
      node1584 = node1580_r;
      node1585_r = node1571_r & pixel[439];
      node1585_l = node1571_r & ~pixel[439];
      node1586_r = node1585_l & pixel[413];
      node1586_l = node1585_l & ~pixel[413];
      node1587 = node1586_l;
      node1588 = node1586_r;
      node1589 = node1585_r;
      node1590_r = node1570_r & pixel[299];
      node1590_l = node1570_r & ~pixel[299];
      node1591_r = node1590_l & pixel[104];
      node1591_l = node1590_l & ~pixel[104];
      node1592_r = node1591_l & pixel[316];
      node1592_l = node1591_l & ~pixel[316];
      node1593_r = node1592_l & pixel[604];
      node1593_l = node1592_l & ~pixel[604];
      node1594 = node1593_l;
      node1595 = node1593_r;
      node1596_r = node1592_r & pixel[216];
      node1596_l = node1592_r & ~pixel[216];
      node1597 = node1596_l;
      node1598 = node1596_r;
      node1599 = node1591_r;
      node1600_r = node1590_r & pixel[604];
      node1600_l = node1590_r & ~pixel[604];
      node1601_r = node1600_l & pixel[270];
      node1601_l = node1600_l & ~pixel[270];
      node1602 = node1601_l;
      node1603_r = node1601_r & pixel[344];
      node1603_l = node1601_r & ~pixel[344];
      node1604 = node1603_l;
      node1605 = node1603_r;
      node1606_r = node1600_r & pixel[345];
      node1606_l = node1600_r & ~pixel[345];
      node1607_r = node1606_l & pixel[383];
      node1607_l = node1606_l & ~pixel[383];
      node1608 = node1607_l;
      node1609 = node1607_r;
      node1610_r = node1606_r & pixel[525];
      node1610_l = node1606_r & ~pixel[525];
      node1611 = node1610_l;
      node1612 = node1610_r;
      result0 = node18 | node42 | node54 | node56 | node69 | node73 | node75 | node79 | node85 | node90 | node91 | node93 | node250 | node259 | node263 | node451 | node458 | node461 | node535 | node614 | node645 | node657 | node672 | node693 | node700 | node703 | node751 | node754 | node799 | node813 | node814 | node816 | node817 | node858 | node889 | node892 | node928 | node955 | node985 | node987 | node993 | node994 | node1102 | node1117 | node1126 | node1127 | node1136 | node1149 | node1156 | node1159 | node1162 | node1163 | node1177 | node1208 | node1217 | node1230 | node1236 | node1239 | node1292 | node1315 | node1331 | node1333 | node1362 | node1365 | node1367 | node1375 | node1377 | node1385 | node1388 | node1395 | node1397 | node1419 | node1420 | node1427 | node1428 | node1431 | node1444 | node1446 | node1452 | node1453 | node1454 | node1458 | node1463 | node1464 | node1466 | node1467 | node1470 | node1473 | node1505 | node1531 | node1582 | node1605 | node1608 | node1611 | node1612;
      result1 = node21 | node211 | node214 | node218 | node224 | node225 | node228 | node241 | node255 | node286 | node303 | node355 | node417 | node421 | node904 | node915 | node920 | node1065 | node1080 | node1094 | node1359;
      result2 = node41 | node46 | node101 | node112 | node137 | node158 | node175 | node189 | node212 | node231 | node235 | node240 | node247 | node264 | node363 | node411 | node422 | node438 | node470 | node530 | node531 | node538 | node542 | node545 | node675 | node686 | node706 | node715 | node722 | node725 | node747 | node764 | node897 | node899 | node908 | node911 | node912 | node927 | node935 | node942 | node952 | node959 | node960 | node967 | node968 | node971 | node981 | node1006 | node1013 | node1033 | node1036 | node1052 | node1072 | node1075 | node1076 | node1083 | node1086 | node1088 | node1089 | node1098 | node1105 | node1109 | node1112 | node1113 | node1118 | node1130 | node1141 | node1147 | node1171 | node1201 | node1247 | node1257 | node1261 | node1263 | node1270 | node1271 | node1277 | node1284 | node1291 | node1298 | node1299 | node1301 | node1305 | node1306 | node1309 | node1327 | node1339 | node1342 | node1373 | node1387 | node1389 | node1398 | node1404 | node1408 | node1414 | node1435 | node1471 | node1482 | node1485 | node1503 | node1523 | node1526 | node1530 | node1541 | node1547 | node1563 | node1568 | node1589 | node1594 | node1604;
      result3 = node63 | node66 | node84 | node94 | node243 | node244 | node270 | node274 | node289 | node295 | node296 | node298 | node304 | node308 | node311 | node312 | node315 | node316 | node318 | node343 | node347 | node349 | node350 | node387 | node388 | node397 | node402 | node410 | node413 | node416 | node425 | node439 | node445 | node460 | node466 | node469 | node473 | node476 | node477 | node484 | node514 | node516 | node537 | node543 | node546 | node549 | node568 | node629 | node687 | node828 | node841 | node852 | node854 | node859 | node866 | node872 | node893 | node956 | node962 | node977 | node980 | node1002 | node1003 | node1005 | node1012 | node1025 | node1028 | node1034 | node1037 | node1040 | node1041 | node1044 | node1049 | node1051 | node1059 | node1137 | node1144 | node1158 | node1183 | node1191 | node1198 | node1202 | node1214 | node1218 | node1222 | node1224 | node1233 | node1237 | node1278 | node1308 | node1314 | node1319 | node1330 | node1407 | node1418 | node1493 | node1584;
      result4 = node11 | node20 | node126 | node127 | node136 | node141 | node145 | node152 | node161 | node184 | node185 | node200 | node326 | node426 | node435 | node436 | node450 | node481 | node491 | node501 | node502 | node505 | node506 | node508 | node513 | node529 | node560 | node567 | node570 | node578 | node589 | node594 | node597 | node603 | node607 | node621 | node653 | node656 | node683 | node721 | node732 | node740 | node752 | node763 | node809 | node821 | node875 | node938 | node995 | node1081 | node1084 | node1273 | node1282 | node1322 | node1338 | node1436 | node1514 | node1539 | node1555 | node1564 | node1578;
      result5 = node17 | node25 | node31 | node49 | node57 | node64 | node67 | node70 | node76 | node86 | node89 | node102 | node149 | node162 | node174 | node177 | node187 | node194 | node202 | node215 | node219 | node220 | node256 | node262 | node271 | node273 | node282 | node302 | node319 | node334 | node346 | node390 | node394 | node395 | node398 | node403 | node446 | node454 | node457 | node474 | node485 | node488 | node489 | node534 | node550 | node552 | node563 | node571 | node575 | node576 | node583 | node610 | node613 | node618 | node622 | node625 | node635 | node642 | node644 | node736 | node739 | node745 | node768 | node770 | node784 | node787 | node791 | node796 | node802 | node808 | node824 | node842 | node844 | node855 | node865 | node878 | node890 | node896 | node900 | node905 | node930 | node936 | node945 | node963 | node984 | node992 | node1009 | node1010 | node1017 | node1018 | node1020 | node1021 | node1024 | node1043 | node1048 | node1055 | node1058 | node1095 | node1129 | node1133 | node1142 | node1150 | node1168 | node1172 | node1184 | node1186 | node1190 | node1193 | node1194 | node1205 | node1215 | node1229 | node1232 | node1265 | node1288 | node1358 | node1368 | node1379 | node1439 | node1442 | node1459 | node1474 | node1492 | node1497 | node1506;
      result6 = node13 | node14 | node24 | node26 | node38 | node103 | node106 | node107 | node120 | node121 | node129 | node133 | node134 | node178 | node232 | node248 | node251 | node275 | node333 | node335 | node366 | node380 | node453 | node467 | node561 | node590 | node591 | node592 | node596 | node668 | node669 | node671 | node676 | node679 | node699 | node707 | node717 | node718 | node730 | node733 | node737 | node744 | node800 | node939 | node953 | node970 | node972 | node1068 | node1134 | node1155 | node1164 | node1169 | node1174 | node1187 | node1199 | node1248 | node1250 | node1254 | node1255 | node1258 | node1274 | node1279 | node1289 | node1302 | node1341 | node1366 | node1374 | node1396 | node1400 | node1434 | node1441 | node1447 | node1457 | node1475 | node1481 | node1490 | node1538 | node1548 | node1549 | node1559 | node1575 | node1576 | node1579 | node1588 | node1595 | node1597 | node1598 | node1599 | node1602;
      result7 = node10 | node32 | node34 | node35 | node47 | node78 | node113 | node115 | node144 | node159 | node165 | node168 | node169 | node183 | node190 | node279 | node327 | node329 | node342 | node362 | node371 | node423 | node443 | node517 | node579 | node650 | node678 | node775 | node778 | node794 | node861 | node871 | node876 | node924 | node1348 | node1349 | node1380 | node1415 | node1484 | node1489 | node1518;
      result8 = node50 | node108 | node116 | node173 | node195 | node197 | node198 | node203 | node227 | node234 | node258 | node287 | node290 | node299 | node309 | node340 | node356 | node358 | node365 | node370 | node373 | node374 | node381 | node391 | node405 | node521 | node553 | node564 | node581 | node626 | node638 | node660 | node694 | node709 | node710 | node714 | node724 | node748 | node755 | node761 | node767 | node771 | node786 | node790 | node793 | node803 | node810 | node822 | node831 | node832 | node838 | node839 | node846 | node847 | node851 | node862 | node879 | node907 | node914 | node921 | node923 | node931 | node943 | node946 | node978 | node988 | node1027 | node1056 | node1066 | node1069 | node1073 | node1097 | node1101 | node1104 | node1110 | node1115 | node1176 | node1206 | node1209 | node1221 | node1225 | node1251 | node1285 | node1318 | node1321 | node1328 | node1345 | node1346 | node1361 | node1384 | node1401 | node1409 | node1412 | node1430 | node1498 | node1501 | node1512 | node1513 | node1515 | node1521 | node1525 | node1528 | node1542 | node1543 | node1556 | node1557 | node1560 | node1567 | node1569 | node1587;
      result9 = node39 | node53 | node119 | node130 | node142 | node148 | node151 | node166 | node280 | node283 | node330 | node339 | node359 | node377 | node378 | node404 | node414 | node442 | node482 | node492 | node498 | node499 | node509 | node520 | node523 | node524 | node584 | node604 | node606 | node611 | node619 | node628 | node634 | node637 | node641 | node649 | node652 | node659 | node684 | node690 | node691 | node702 | node760 | node776 | node777 | node825 | node829 | node869 | node1145 | node1240 | node1264 | node1312 | node1334 | node1500 | node1517 | node1550 | node1583 | node1609;

      tree_1 = {result9, result8, result7, result6, result5, result4, result3, result2, result1, result0};
    end
  endfunction

  function [9:0] tree_2;
    input [783:0] pixel;

    reg node0_r;
    reg node0_l;
    reg node1_r;
    reg node1_l;
    reg node2_r;
    reg node2_l;
    reg node3_r;
    reg node3_l;
    reg node4_r;
    reg node4_l;
    reg node5_r;
    reg node5_l;
    reg node6_r;
    reg node6_l;
    reg node7_r;
    reg node7_l;
    reg node8_r;
    reg node8_l;
    reg node9_r;
    reg node9_l;
    reg node10;
    reg node11;
    reg node12_r;
    reg node12_l;
    reg node13;
    reg node14;
    reg node15_r;
    reg node15_l;
    reg node16_r;
    reg node16_l;
    reg node17;
    reg node18;
    reg node19_r;
    reg node19_l;
    reg node20;
    reg node21;
    reg node22_r;
    reg node22_l;
    reg node23_r;
    reg node23_l;
    reg node24_r;
    reg node24_l;
    reg node25;
    reg node26;
    reg node27_r;
    reg node27_l;
    reg node28;
    reg node29;
    reg node30_r;
    reg node30_l;
    reg node31_r;
    reg node31_l;
    reg node32;
    reg node33;
    reg node34_r;
    reg node34_l;
    reg node35;
    reg node36;
    reg node37_r;
    reg node37_l;
    reg node38_r;
    reg node38_l;
    reg node39_r;
    reg node39_l;
    reg node40_r;
    reg node40_l;
    reg node41;
    reg node42;
    reg node43_r;
    reg node43_l;
    reg node44;
    reg node45;
    reg node46_r;
    reg node46_l;
    reg node47_r;
    reg node47_l;
    reg node48;
    reg node49;
    reg node50_r;
    reg node50_l;
    reg node51;
    reg node52;
    reg node53_r;
    reg node53_l;
    reg node54_r;
    reg node54_l;
    reg node55_r;
    reg node55_l;
    reg node56;
    reg node57;
    reg node58_r;
    reg node58_l;
    reg node59;
    reg node60;
    reg node61_r;
    reg node61_l;
    reg node62_r;
    reg node62_l;
    reg node63;
    reg node64;
    reg node65_r;
    reg node65_l;
    reg node66;
    reg node67;
    reg node68_r;
    reg node68_l;
    reg node69_r;
    reg node69_l;
    reg node70_r;
    reg node70_l;
    reg node71_r;
    reg node71_l;
    reg node72_r;
    reg node72_l;
    reg node73;
    reg node74;
    reg node75_r;
    reg node75_l;
    reg node76;
    reg node77;
    reg node78_r;
    reg node78_l;
    reg node79_r;
    reg node79_l;
    reg node80;
    reg node81;
    reg node82_r;
    reg node82_l;
    reg node83;
    reg node84;
    reg node85_r;
    reg node85_l;
    reg node86_r;
    reg node86_l;
    reg node87_r;
    reg node87_l;
    reg node88;
    reg node89;
    reg node90_r;
    reg node90_l;
    reg node91;
    reg node92;
    reg node93_r;
    reg node93_l;
    reg node94_r;
    reg node94_l;
    reg node95;
    reg node96;
    reg node97_r;
    reg node97_l;
    reg node98;
    reg node99;
    reg node100_r;
    reg node100_l;
    reg node101_r;
    reg node101_l;
    reg node102;
    reg node103_r;
    reg node103_l;
    reg node104_r;
    reg node104_l;
    reg node105;
    reg node106;
    reg node107;
    reg node108_r;
    reg node108_l;
    reg node109;
    reg node110_r;
    reg node110_l;
    reg node111;
    reg node112;
    reg node113_r;
    reg node113_l;
    reg node114_r;
    reg node114_l;
    reg node115_r;
    reg node115_l;
    reg node116_r;
    reg node116_l;
    reg node117_r;
    reg node117_l;
    reg node118_r;
    reg node118_l;
    reg node119;
    reg node120;
    reg node121_r;
    reg node121_l;
    reg node122;
    reg node123;
    reg node124_r;
    reg node124_l;
    reg node125_r;
    reg node125_l;
    reg node126;
    reg node127;
    reg node128_r;
    reg node128_l;
    reg node129;
    reg node130;
    reg node131_r;
    reg node131_l;
    reg node132_r;
    reg node132_l;
    reg node133_r;
    reg node133_l;
    reg node134;
    reg node135;
    reg node136_r;
    reg node136_l;
    reg node137;
    reg node138;
    reg node139_r;
    reg node139_l;
    reg node140_r;
    reg node140_l;
    reg node141;
    reg node142;
    reg node143_r;
    reg node143_l;
    reg node144;
    reg node145;
    reg node146_r;
    reg node146_l;
    reg node147_r;
    reg node147_l;
    reg node148_r;
    reg node148_l;
    reg node149_r;
    reg node149_l;
    reg node150;
    reg node151;
    reg node152_r;
    reg node152_l;
    reg node153;
    reg node154;
    reg node155_r;
    reg node155_l;
    reg node156_r;
    reg node156_l;
    reg node157;
    reg node158;
    reg node159;
    reg node160_r;
    reg node160_l;
    reg node161_r;
    reg node161_l;
    reg node162_r;
    reg node162_l;
    reg node163;
    reg node164;
    reg node165_r;
    reg node165_l;
    reg node166;
    reg node167;
    reg node168_r;
    reg node168_l;
    reg node169_r;
    reg node169_l;
    reg node170;
    reg node171;
    reg node172_r;
    reg node172_l;
    reg node173;
    reg node174;
    reg node175_r;
    reg node175_l;
    reg node176_r;
    reg node176_l;
    reg node177_r;
    reg node177_l;
    reg node178_r;
    reg node178_l;
    reg node179_r;
    reg node179_l;
    reg node180;
    reg node181;
    reg node182_r;
    reg node182_l;
    reg node183;
    reg node184;
    reg node185_r;
    reg node185_l;
    reg node186_r;
    reg node186_l;
    reg node187;
    reg node188;
    reg node189;
    reg node190_r;
    reg node190_l;
    reg node191_r;
    reg node191_l;
    reg node192_r;
    reg node192_l;
    reg node193;
    reg node194;
    reg node195_r;
    reg node195_l;
    reg node196;
    reg node197;
    reg node198_r;
    reg node198_l;
    reg node199_r;
    reg node199_l;
    reg node200;
    reg node201;
    reg node202_r;
    reg node202_l;
    reg node203;
    reg node204;
    reg node205_r;
    reg node205_l;
    reg node206_r;
    reg node206_l;
    reg node207_r;
    reg node207_l;
    reg node208;
    reg node209_r;
    reg node209_l;
    reg node210;
    reg node211;
    reg node212;
    reg node213_r;
    reg node213_l;
    reg node214_r;
    reg node214_l;
    reg node215_r;
    reg node215_l;
    reg node216;
    reg node217;
    reg node218_r;
    reg node218_l;
    reg node219;
    reg node220;
    reg node221;
    reg node222_r;
    reg node222_l;
    reg node223_r;
    reg node223_l;
    reg node224_r;
    reg node224_l;
    reg node225_r;
    reg node225_l;
    reg node226_r;
    reg node226_l;
    reg node227_r;
    reg node227_l;
    reg node228_r;
    reg node228_l;
    reg node229;
    reg node230;
    reg node231_r;
    reg node231_l;
    reg node232;
    reg node233;
    reg node234_r;
    reg node234_l;
    reg node235_r;
    reg node235_l;
    reg node236;
    reg node237;
    reg node238_r;
    reg node238_l;
    reg node239;
    reg node240;
    reg node241_r;
    reg node241_l;
    reg node242_r;
    reg node242_l;
    reg node243_r;
    reg node243_l;
    reg node244;
    reg node245;
    reg node246_r;
    reg node246_l;
    reg node247;
    reg node248;
    reg node249_r;
    reg node249_l;
    reg node250_r;
    reg node250_l;
    reg node251;
    reg node252;
    reg node253_r;
    reg node253_l;
    reg node254;
    reg node255;
    reg node256_r;
    reg node256_l;
    reg node257_r;
    reg node257_l;
    reg node258_r;
    reg node258_l;
    reg node259_r;
    reg node259_l;
    reg node260;
    reg node261;
    reg node262;
    reg node263_r;
    reg node263_l;
    reg node264_r;
    reg node264_l;
    reg node265;
    reg node266;
    reg node267_r;
    reg node267_l;
    reg node268;
    reg node269;
    reg node270_r;
    reg node270_l;
    reg node271_r;
    reg node271_l;
    reg node272_r;
    reg node272_l;
    reg node273;
    reg node274;
    reg node275_r;
    reg node275_l;
    reg node276;
    reg node277;
    reg node278_r;
    reg node278_l;
    reg node279_r;
    reg node279_l;
    reg node280;
    reg node281;
    reg node282_r;
    reg node282_l;
    reg node283;
    reg node284;
    reg node285_r;
    reg node285_l;
    reg node286_r;
    reg node286_l;
    reg node287_r;
    reg node287_l;
    reg node288_r;
    reg node288_l;
    reg node289_r;
    reg node289_l;
    reg node290;
    reg node291;
    reg node292_r;
    reg node292_l;
    reg node293;
    reg node294;
    reg node295_r;
    reg node295_l;
    reg node296_r;
    reg node296_l;
    reg node297;
    reg node298;
    reg node299_r;
    reg node299_l;
    reg node300;
    reg node301;
    reg node302_r;
    reg node302_l;
    reg node303_r;
    reg node303_l;
    reg node304_r;
    reg node304_l;
    reg node305;
    reg node306;
    reg node307_r;
    reg node307_l;
    reg node308;
    reg node309;
    reg node310_r;
    reg node310_l;
    reg node311_r;
    reg node311_l;
    reg node312;
    reg node313;
    reg node314_r;
    reg node314_l;
    reg node315;
    reg node316;
    reg node317_r;
    reg node317_l;
    reg node318_r;
    reg node318_l;
    reg node319_r;
    reg node319_l;
    reg node320;
    reg node321_r;
    reg node321_l;
    reg node322;
    reg node323;
    reg node324_r;
    reg node324_l;
    reg node325;
    reg node326;
    reg node327_r;
    reg node327_l;
    reg node328_r;
    reg node328_l;
    reg node329_r;
    reg node329_l;
    reg node330;
    reg node331;
    reg node332_r;
    reg node332_l;
    reg node333;
    reg node334;
    reg node335;
    reg node336_r;
    reg node336_l;
    reg node337_r;
    reg node337_l;
    reg node338_r;
    reg node338_l;
    reg node339_r;
    reg node339_l;
    reg node340_r;
    reg node340_l;
    reg node341_r;
    reg node341_l;
    reg node342;
    reg node343;
    reg node344;
    reg node345_r;
    reg node345_l;
    reg node346_r;
    reg node346_l;
    reg node347;
    reg node348;
    reg node349_r;
    reg node349_l;
    reg node350;
    reg node351;
    reg node352_r;
    reg node352_l;
    reg node353_r;
    reg node353_l;
    reg node354_r;
    reg node354_l;
    reg node355;
    reg node356;
    reg node357_r;
    reg node357_l;
    reg node358;
    reg node359;
    reg node360_r;
    reg node360_l;
    reg node361_r;
    reg node361_l;
    reg node362;
    reg node363;
    reg node364;
    reg node365_r;
    reg node365_l;
    reg node366_r;
    reg node366_l;
    reg node367_r;
    reg node367_l;
    reg node368;
    reg node369_r;
    reg node369_l;
    reg node370;
    reg node371;
    reg node372_r;
    reg node372_l;
    reg node373_r;
    reg node373_l;
    reg node374;
    reg node375;
    reg node376_r;
    reg node376_l;
    reg node377;
    reg node378;
    reg node379_r;
    reg node379_l;
    reg node380_r;
    reg node380_l;
    reg node381_r;
    reg node381_l;
    reg node382;
    reg node383;
    reg node384_r;
    reg node384_l;
    reg node385;
    reg node386;
    reg node387_r;
    reg node387_l;
    reg node388_r;
    reg node388_l;
    reg node389;
    reg node390;
    reg node391_r;
    reg node391_l;
    reg node392;
    reg node393;
    reg node394_r;
    reg node394_l;
    reg node395_r;
    reg node395_l;
    reg node396_r;
    reg node396_l;
    reg node397_r;
    reg node397_l;
    reg node398_r;
    reg node398_l;
    reg node399;
    reg node400;
    reg node401_r;
    reg node401_l;
    reg node402;
    reg node403;
    reg node404_r;
    reg node404_l;
    reg node405_r;
    reg node405_l;
    reg node406;
    reg node407;
    reg node408_r;
    reg node408_l;
    reg node409;
    reg node410;
    reg node411_r;
    reg node411_l;
    reg node412;
    reg node413_r;
    reg node413_l;
    reg node414_r;
    reg node414_l;
    reg node415;
    reg node416;
    reg node417;
    reg node418_r;
    reg node418_l;
    reg node419_r;
    reg node419_l;
    reg node420_r;
    reg node420_l;
    reg node421_r;
    reg node421_l;
    reg node422;
    reg node423;
    reg node424_r;
    reg node424_l;
    reg node425;
    reg node426;
    reg node427_r;
    reg node427_l;
    reg node428_r;
    reg node428_l;
    reg node429;
    reg node430;
    reg node431_r;
    reg node431_l;
    reg node432;
    reg node433;
    reg node434_r;
    reg node434_l;
    reg node435_r;
    reg node435_l;
    reg node436_r;
    reg node436_l;
    reg node437;
    reg node438;
    reg node439_r;
    reg node439_l;
    reg node440;
    reg node441;
    reg node442_r;
    reg node442_l;
    reg node443_r;
    reg node443_l;
    reg node444;
    reg node445;
    reg node446_r;
    reg node446_l;
    reg node447;
    reg node448;
    reg node449_r;
    reg node449_l;
    reg node450_r;
    reg node450_l;
    reg node451_r;
    reg node451_l;
    reg node452_r;
    reg node452_l;
    reg node453_r;
    reg node453_l;
    reg node454_r;
    reg node454_l;
    reg node455_r;
    reg node455_l;
    reg node456_r;
    reg node456_l;
    reg node457;
    reg node458;
    reg node459_r;
    reg node459_l;
    reg node460;
    reg node461;
    reg node462_r;
    reg node462_l;
    reg node463_r;
    reg node463_l;
    reg node464;
    reg node465;
    reg node466_r;
    reg node466_l;
    reg node467;
    reg node468;
    reg node469_r;
    reg node469_l;
    reg node470_r;
    reg node470_l;
    reg node471;
    reg node472;
    reg node473;
    reg node474_r;
    reg node474_l;
    reg node475_r;
    reg node475_l;
    reg node476_r;
    reg node476_l;
    reg node477_r;
    reg node477_l;
    reg node478;
    reg node479;
    reg node480_r;
    reg node480_l;
    reg node481;
    reg node482;
    reg node483_r;
    reg node483_l;
    reg node484_r;
    reg node484_l;
    reg node485;
    reg node486;
    reg node487_r;
    reg node487_l;
    reg node488;
    reg node489;
    reg node490_r;
    reg node490_l;
    reg node491_r;
    reg node491_l;
    reg node492_r;
    reg node492_l;
    reg node493;
    reg node494;
    reg node495;
    reg node496;
    reg node497_r;
    reg node497_l;
    reg node498_r;
    reg node498_l;
    reg node499_r;
    reg node499_l;
    reg node500_r;
    reg node500_l;
    reg node501_r;
    reg node501_l;
    reg node502;
    reg node503;
    reg node504_r;
    reg node504_l;
    reg node505;
    reg node506;
    reg node507_r;
    reg node507_l;
    reg node508_r;
    reg node508_l;
    reg node509;
    reg node510;
    reg node511;
    reg node512_r;
    reg node512_l;
    reg node513_r;
    reg node513_l;
    reg node514_r;
    reg node514_l;
    reg node515;
    reg node516;
    reg node517_r;
    reg node517_l;
    reg node518;
    reg node519;
    reg node520_r;
    reg node520_l;
    reg node521_r;
    reg node521_l;
    reg node522;
    reg node523;
    reg node524;
    reg node525_r;
    reg node525_l;
    reg node526_r;
    reg node526_l;
    reg node527_r;
    reg node527_l;
    reg node528_r;
    reg node528_l;
    reg node529;
    reg node530;
    reg node531;
    reg node532;
    reg node533;
    reg node534_r;
    reg node534_l;
    reg node535_r;
    reg node535_l;
    reg node536_r;
    reg node536_l;
    reg node537_r;
    reg node537_l;
    reg node538_r;
    reg node538_l;
    reg node539_r;
    reg node539_l;
    reg node540;
    reg node541;
    reg node542_r;
    reg node542_l;
    reg node543;
    reg node544;
    reg node545_r;
    reg node545_l;
    reg node546;
    reg node547_r;
    reg node547_l;
    reg node548;
    reg node549;
    reg node550_r;
    reg node550_l;
    reg node551_r;
    reg node551_l;
    reg node552_r;
    reg node552_l;
    reg node553;
    reg node554;
    reg node555_r;
    reg node555_l;
    reg node556;
    reg node557;
    reg node558_r;
    reg node558_l;
    reg node559_r;
    reg node559_l;
    reg node560;
    reg node561;
    reg node562;
    reg node563_r;
    reg node563_l;
    reg node564_r;
    reg node564_l;
    reg node565_r;
    reg node565_l;
    reg node566_r;
    reg node566_l;
    reg node567;
    reg node568;
    reg node569_r;
    reg node569_l;
    reg node570;
    reg node571;
    reg node572_r;
    reg node572_l;
    reg node573_r;
    reg node573_l;
    reg node574;
    reg node575;
    reg node576_r;
    reg node576_l;
    reg node577;
    reg node578;
    reg node579_r;
    reg node579_l;
    reg node580_r;
    reg node580_l;
    reg node581_r;
    reg node581_l;
    reg node582;
    reg node583;
    reg node584_r;
    reg node584_l;
    reg node585;
    reg node586;
    reg node587_r;
    reg node587_l;
    reg node588_r;
    reg node588_l;
    reg node589;
    reg node590;
    reg node591_r;
    reg node591_l;
    reg node592;
    reg node593;
    reg node594_r;
    reg node594_l;
    reg node595_r;
    reg node595_l;
    reg node596_r;
    reg node596_l;
    reg node597_r;
    reg node597_l;
    reg node598_r;
    reg node598_l;
    reg node599;
    reg node600;
    reg node601;
    reg node602_r;
    reg node602_l;
    reg node603_r;
    reg node603_l;
    reg node604;
    reg node605;
    reg node606_r;
    reg node606_l;
    reg node607;
    reg node608;
    reg node609_r;
    reg node609_l;
    reg node610_r;
    reg node610_l;
    reg node611_r;
    reg node611_l;
    reg node612;
    reg node613;
    reg node614_r;
    reg node614_l;
    reg node615;
    reg node616;
    reg node617_r;
    reg node617_l;
    reg node618_r;
    reg node618_l;
    reg node619;
    reg node620;
    reg node621_r;
    reg node621_l;
    reg node622;
    reg node623;
    reg node624_r;
    reg node624_l;
    reg node625;
    reg node626_r;
    reg node626_l;
    reg node627;
    reg node628_r;
    reg node628_l;
    reg node629_r;
    reg node629_l;
    reg node630;
    reg node631;
    reg node632;
    reg node633_r;
    reg node633_l;
    reg node634_r;
    reg node634_l;
    reg node635_r;
    reg node635_l;
    reg node636_r;
    reg node636_l;
    reg node637_r;
    reg node637_l;
    reg node638_r;
    reg node638_l;
    reg node639_r;
    reg node639_l;
    reg node640;
    reg node641;
    reg node642_r;
    reg node642_l;
    reg node643;
    reg node644;
    reg node645_r;
    reg node645_l;
    reg node646_r;
    reg node646_l;
    reg node647;
    reg node648;
    reg node649_r;
    reg node649_l;
    reg node650;
    reg node651;
    reg node652_r;
    reg node652_l;
    reg node653_r;
    reg node653_l;
    reg node654_r;
    reg node654_l;
    reg node655;
    reg node656;
    reg node657_r;
    reg node657_l;
    reg node658;
    reg node659;
    reg node660_r;
    reg node660_l;
    reg node661_r;
    reg node661_l;
    reg node662;
    reg node663;
    reg node664_r;
    reg node664_l;
    reg node665;
    reg node666;
    reg node667_r;
    reg node667_l;
    reg node668_r;
    reg node668_l;
    reg node669_r;
    reg node669_l;
    reg node670_r;
    reg node670_l;
    reg node671;
    reg node672;
    reg node673_r;
    reg node673_l;
    reg node674;
    reg node675;
    reg node676_r;
    reg node676_l;
    reg node677_r;
    reg node677_l;
    reg node678;
    reg node679;
    reg node680;
    reg node681_r;
    reg node681_l;
    reg node682_r;
    reg node682_l;
    reg node683_r;
    reg node683_l;
    reg node684;
    reg node685;
    reg node686_r;
    reg node686_l;
    reg node687;
    reg node688;
    reg node689_r;
    reg node689_l;
    reg node690_r;
    reg node690_l;
    reg node691;
    reg node692;
    reg node693_r;
    reg node693_l;
    reg node694;
    reg node695;
    reg node696_r;
    reg node696_l;
    reg node697_r;
    reg node697_l;
    reg node698_r;
    reg node698_l;
    reg node699_r;
    reg node699_l;
    reg node700_r;
    reg node700_l;
    reg node701;
    reg node702;
    reg node703_r;
    reg node703_l;
    reg node704;
    reg node705;
    reg node706_r;
    reg node706_l;
    reg node707_r;
    reg node707_l;
    reg node708;
    reg node709;
    reg node710_r;
    reg node710_l;
    reg node711;
    reg node712;
    reg node713_r;
    reg node713_l;
    reg node714_r;
    reg node714_l;
    reg node715_r;
    reg node715_l;
    reg node716;
    reg node717;
    reg node718_r;
    reg node718_l;
    reg node719;
    reg node720;
    reg node721_r;
    reg node721_l;
    reg node722_r;
    reg node722_l;
    reg node723;
    reg node724;
    reg node725_r;
    reg node725_l;
    reg node726;
    reg node727;
    reg node728_r;
    reg node728_l;
    reg node729_r;
    reg node729_l;
    reg node730_r;
    reg node730_l;
    reg node731_r;
    reg node731_l;
    reg node732;
    reg node733;
    reg node734_r;
    reg node734_l;
    reg node735;
    reg node736;
    reg node737_r;
    reg node737_l;
    reg node738;
    reg node739_r;
    reg node739_l;
    reg node740;
    reg node741;
    reg node742_r;
    reg node742_l;
    reg node743_r;
    reg node743_l;
    reg node744_r;
    reg node744_l;
    reg node745;
    reg node746;
    reg node747_r;
    reg node747_l;
    reg node748;
    reg node749;
    reg node750;
    reg node751_r;
    reg node751_l;
    reg node752_r;
    reg node752_l;
    reg node753_r;
    reg node753_l;
    reg node754_r;
    reg node754_l;
    reg node755_r;
    reg node755_l;
    reg node756_r;
    reg node756_l;
    reg node757;
    reg node758;
    reg node759_r;
    reg node759_l;
    reg node760;
    reg node761;
    reg node762_r;
    reg node762_l;
    reg node763_r;
    reg node763_l;
    reg node764;
    reg node765;
    reg node766_r;
    reg node766_l;
    reg node767;
    reg node768;
    reg node769_r;
    reg node769_l;
    reg node770_r;
    reg node770_l;
    reg node771_r;
    reg node771_l;
    reg node772;
    reg node773;
    reg node774_r;
    reg node774_l;
    reg node775;
    reg node776;
    reg node777_r;
    reg node777_l;
    reg node778_r;
    reg node778_l;
    reg node779;
    reg node780;
    reg node781_r;
    reg node781_l;
    reg node782;
    reg node783;
    reg node784_r;
    reg node784_l;
    reg node785_r;
    reg node785_l;
    reg node786_r;
    reg node786_l;
    reg node787_r;
    reg node787_l;
    reg node788;
    reg node789;
    reg node790_r;
    reg node790_l;
    reg node791;
    reg node792;
    reg node793_r;
    reg node793_l;
    reg node794_r;
    reg node794_l;
    reg node795;
    reg node796;
    reg node797_r;
    reg node797_l;
    reg node798;
    reg node799;
    reg node800_r;
    reg node800_l;
    reg node801_r;
    reg node801_l;
    reg node802_r;
    reg node802_l;
    reg node803;
    reg node804;
    reg node805_r;
    reg node805_l;
    reg node806;
    reg node807;
    reg node808_r;
    reg node808_l;
    reg node809;
    reg node810_r;
    reg node810_l;
    reg node811;
    reg node812;
    reg node813_r;
    reg node813_l;
    reg node814_r;
    reg node814_l;
    reg node815_r;
    reg node815_l;
    reg node816_r;
    reg node816_l;
    reg node817_r;
    reg node817_l;
    reg node818;
    reg node819;
    reg node820_r;
    reg node820_l;
    reg node821;
    reg node822;
    reg node823_r;
    reg node823_l;
    reg node824_r;
    reg node824_l;
    reg node825;
    reg node826;
    reg node827_r;
    reg node827_l;
    reg node828;
    reg node829;
    reg node830_r;
    reg node830_l;
    reg node831_r;
    reg node831_l;
    reg node832_r;
    reg node832_l;
    reg node833;
    reg node834;
    reg node835_r;
    reg node835_l;
    reg node836;
    reg node837;
    reg node838_r;
    reg node838_l;
    reg node839_r;
    reg node839_l;
    reg node840;
    reg node841;
    reg node842_r;
    reg node842_l;
    reg node843;
    reg node844;
    reg node845_r;
    reg node845_l;
    reg node846_r;
    reg node846_l;
    reg node847_r;
    reg node847_l;
    reg node848_r;
    reg node848_l;
    reg node849;
    reg node850;
    reg node851_r;
    reg node851_l;
    reg node852;
    reg node853;
    reg node854_r;
    reg node854_l;
    reg node855_r;
    reg node855_l;
    reg node856;
    reg node857;
    reg node858_r;
    reg node858_l;
    reg node859;
    reg node860;
    reg node861_r;
    reg node861_l;
    reg node862_r;
    reg node862_l;
    reg node863_r;
    reg node863_l;
    reg node864;
    reg node865;
    reg node866_r;
    reg node866_l;
    reg node867;
    reg node868;
    reg node869_r;
    reg node869_l;
    reg node870_r;
    reg node870_l;
    reg node871;
    reg node872;
    reg node873_r;
    reg node873_l;
    reg node874;
    reg node875;
    reg node876_r;
    reg node876_l;
    reg node877_r;
    reg node877_l;
    reg node878_r;
    reg node878_l;
    reg node879_r;
    reg node879_l;
    reg node880_r;
    reg node880_l;
    reg node881_r;
    reg node881_l;
    reg node882_r;
    reg node882_l;
    reg node883_r;
    reg node883_l;
    reg node884_r;
    reg node884_l;
    reg node885;
    reg node886;
    reg node887_r;
    reg node887_l;
    reg node888;
    reg node889;
    reg node890_r;
    reg node890_l;
    reg node891_r;
    reg node891_l;
    reg node892;
    reg node893;
    reg node894_r;
    reg node894_l;
    reg node895;
    reg node896;
    reg node897_r;
    reg node897_l;
    reg node898_r;
    reg node898_l;
    reg node899_r;
    reg node899_l;
    reg node900;
    reg node901;
    reg node902_r;
    reg node902_l;
    reg node903;
    reg node904;
    reg node905_r;
    reg node905_l;
    reg node906_r;
    reg node906_l;
    reg node907;
    reg node908;
    reg node909_r;
    reg node909_l;
    reg node910;
    reg node911;
    reg node912_r;
    reg node912_l;
    reg node913_r;
    reg node913_l;
    reg node914_r;
    reg node914_l;
    reg node915_r;
    reg node915_l;
    reg node916;
    reg node917;
    reg node918_r;
    reg node918_l;
    reg node919;
    reg node920;
    reg node921_r;
    reg node921_l;
    reg node922_r;
    reg node922_l;
    reg node923;
    reg node924;
    reg node925_r;
    reg node925_l;
    reg node926;
    reg node927;
    reg node928_r;
    reg node928_l;
    reg node929_r;
    reg node929_l;
    reg node930;
    reg node931_r;
    reg node931_l;
    reg node932;
    reg node933;
    reg node934_r;
    reg node934_l;
    reg node935_r;
    reg node935_l;
    reg node936;
    reg node937;
    reg node938_r;
    reg node938_l;
    reg node939;
    reg node940;
    reg node941_r;
    reg node941_l;
    reg node942_r;
    reg node942_l;
    reg node943_r;
    reg node943_l;
    reg node944_r;
    reg node944_l;
    reg node945_r;
    reg node945_l;
    reg node946;
    reg node947;
    reg node948_r;
    reg node948_l;
    reg node949;
    reg node950;
    reg node951_r;
    reg node951_l;
    reg node952_r;
    reg node952_l;
    reg node953;
    reg node954;
    reg node955_r;
    reg node955_l;
    reg node956;
    reg node957;
    reg node958_r;
    reg node958_l;
    reg node959_r;
    reg node959_l;
    reg node960_r;
    reg node960_l;
    reg node961;
    reg node962;
    reg node963_r;
    reg node963_l;
    reg node964;
    reg node965;
    reg node966_r;
    reg node966_l;
    reg node967_r;
    reg node967_l;
    reg node968;
    reg node969;
    reg node970_r;
    reg node970_l;
    reg node971;
    reg node972;
    reg node973_r;
    reg node973_l;
    reg node974_r;
    reg node974_l;
    reg node975_r;
    reg node975_l;
    reg node976_r;
    reg node976_l;
    reg node977;
    reg node978;
    reg node979_r;
    reg node979_l;
    reg node980;
    reg node981;
    reg node982_r;
    reg node982_l;
    reg node983_r;
    reg node983_l;
    reg node984;
    reg node985;
    reg node986_r;
    reg node986_l;
    reg node987;
    reg node988;
    reg node989_r;
    reg node989_l;
    reg node990_r;
    reg node990_l;
    reg node991_r;
    reg node991_l;
    reg node992;
    reg node993;
    reg node994;
    reg node995_r;
    reg node995_l;
    reg node996;
    reg node997_r;
    reg node997_l;
    reg node998;
    reg node999;
    reg node1000_r;
    reg node1000_l;
    reg node1001_r;
    reg node1001_l;
    reg node1002_r;
    reg node1002_l;
    reg node1003_r;
    reg node1003_l;
    reg node1004_r;
    reg node1004_l;
    reg node1005_r;
    reg node1005_l;
    reg node1006;
    reg node1007;
    reg node1008_r;
    reg node1008_l;
    reg node1009;
    reg node1010;
    reg node1011_r;
    reg node1011_l;
    reg node1012_r;
    reg node1012_l;
    reg node1013;
    reg node1014;
    reg node1015_r;
    reg node1015_l;
    reg node1016;
    reg node1017;
    reg node1018_r;
    reg node1018_l;
    reg node1019_r;
    reg node1019_l;
    reg node1020_r;
    reg node1020_l;
    reg node1021;
    reg node1022;
    reg node1023_r;
    reg node1023_l;
    reg node1024;
    reg node1025;
    reg node1026_r;
    reg node1026_l;
    reg node1027;
    reg node1028;
    reg node1029_r;
    reg node1029_l;
    reg node1030_r;
    reg node1030_l;
    reg node1031_r;
    reg node1031_l;
    reg node1032_r;
    reg node1032_l;
    reg node1033;
    reg node1034;
    reg node1035_r;
    reg node1035_l;
    reg node1036;
    reg node1037;
    reg node1038_r;
    reg node1038_l;
    reg node1039_r;
    reg node1039_l;
    reg node1040;
    reg node1041;
    reg node1042;
    reg node1043_r;
    reg node1043_l;
    reg node1044_r;
    reg node1044_l;
    reg node1045_r;
    reg node1045_l;
    reg node1046;
    reg node1047;
    reg node1048_r;
    reg node1048_l;
    reg node1049;
    reg node1050;
    reg node1051_r;
    reg node1051_l;
    reg node1052;
    reg node1053;
    reg node1054_r;
    reg node1054_l;
    reg node1055_r;
    reg node1055_l;
    reg node1056_r;
    reg node1056_l;
    reg node1057_r;
    reg node1057_l;
    reg node1058_r;
    reg node1058_l;
    reg node1059;
    reg node1060;
    reg node1061;
    reg node1062;
    reg node1063_r;
    reg node1063_l;
    reg node1064_r;
    reg node1064_l;
    reg node1065;
    reg node1066_r;
    reg node1066_l;
    reg node1067;
    reg node1068;
    reg node1069_r;
    reg node1069_l;
    reg node1070_r;
    reg node1070_l;
    reg node1071;
    reg node1072;
    reg node1073;
    reg node1074_r;
    reg node1074_l;
    reg node1075_r;
    reg node1075_l;
    reg node1076_r;
    reg node1076_l;
    reg node1077_r;
    reg node1077_l;
    reg node1078;
    reg node1079;
    reg node1080_r;
    reg node1080_l;
    reg node1081;
    reg node1082;
    reg node1083;
    reg node1084_r;
    reg node1084_l;
    reg node1085_r;
    reg node1085_l;
    reg node1086_r;
    reg node1086_l;
    reg node1087;
    reg node1088;
    reg node1089;
    reg node1090_r;
    reg node1090_l;
    reg node1091_r;
    reg node1091_l;
    reg node1092;
    reg node1093;
    reg node1094;
    reg node1095_r;
    reg node1095_l;
    reg node1096_r;
    reg node1096_l;
    reg node1097_r;
    reg node1097_l;
    reg node1098_r;
    reg node1098_l;
    reg node1099_r;
    reg node1099_l;
    reg node1100_r;
    reg node1100_l;
    reg node1101_r;
    reg node1101_l;
    reg node1102;
    reg node1103;
    reg node1104_r;
    reg node1104_l;
    reg node1105;
    reg node1106;
    reg node1107_r;
    reg node1107_l;
    reg node1108_r;
    reg node1108_l;
    reg node1109;
    reg node1110;
    reg node1111_r;
    reg node1111_l;
    reg node1112;
    reg node1113;
    reg node1114_r;
    reg node1114_l;
    reg node1115_r;
    reg node1115_l;
    reg node1116;
    reg node1117;
    reg node1118;
    reg node1119_r;
    reg node1119_l;
    reg node1120_r;
    reg node1120_l;
    reg node1121_r;
    reg node1121_l;
    reg node1122_r;
    reg node1122_l;
    reg node1123;
    reg node1124;
    reg node1125_r;
    reg node1125_l;
    reg node1126;
    reg node1127;
    reg node1128_r;
    reg node1128_l;
    reg node1129_r;
    reg node1129_l;
    reg node1130;
    reg node1131;
    reg node1132_r;
    reg node1132_l;
    reg node1133;
    reg node1134;
    reg node1135;
    reg node1136_r;
    reg node1136_l;
    reg node1137_r;
    reg node1137_l;
    reg node1138_r;
    reg node1138_l;
    reg node1139_r;
    reg node1139_l;
    reg node1140_r;
    reg node1140_l;
    reg node1141;
    reg node1142;
    reg node1143;
    reg node1144_r;
    reg node1144_l;
    reg node1145_r;
    reg node1145_l;
    reg node1146;
    reg node1147;
    reg node1148;
    reg node1149_r;
    reg node1149_l;
    reg node1150_r;
    reg node1150_l;
    reg node1151_r;
    reg node1151_l;
    reg node1152;
    reg node1153;
    reg node1154_r;
    reg node1154_l;
    reg node1155;
    reg node1156;
    reg node1157;
    reg node1158_r;
    reg node1158_l;
    reg node1159_r;
    reg node1159_l;
    reg node1160_r;
    reg node1160_l;
    reg node1161_r;
    reg node1161_l;
    reg node1162;
    reg node1163;
    reg node1164_r;
    reg node1164_l;
    reg node1165;
    reg node1166;
    reg node1167_r;
    reg node1167_l;
    reg node1168_r;
    reg node1168_l;
    reg node1169;
    reg node1170;
    reg node1171;
    reg node1172_r;
    reg node1172_l;
    reg node1173_r;
    reg node1173_l;
    reg node1174_r;
    reg node1174_l;
    reg node1175;
    reg node1176;
    reg node1177;
    reg node1178_r;
    reg node1178_l;
    reg node1179_r;
    reg node1179_l;
    reg node1180;
    reg node1181;
    reg node1182_r;
    reg node1182_l;
    reg node1183;
    reg node1184;
    reg node1185_r;
    reg node1185_l;
    reg node1186_r;
    reg node1186_l;
    reg node1187_r;
    reg node1187_l;
    reg node1188_r;
    reg node1188_l;
    reg node1189_r;
    reg node1189_l;
    reg node1190_r;
    reg node1190_l;
    reg node1191;
    reg node1192;
    reg node1193_r;
    reg node1193_l;
    reg node1194;
    reg node1195;
    reg node1196_r;
    reg node1196_l;
    reg node1197_r;
    reg node1197_l;
    reg node1198;
    reg node1199;
    reg node1200_r;
    reg node1200_l;
    reg node1201;
    reg node1202;
    reg node1203_r;
    reg node1203_l;
    reg node1204_r;
    reg node1204_l;
    reg node1205_r;
    reg node1205_l;
    reg node1206;
    reg node1207;
    reg node1208;
    reg node1209_r;
    reg node1209_l;
    reg node1210_r;
    reg node1210_l;
    reg node1211;
    reg node1212;
    reg node1213_r;
    reg node1213_l;
    reg node1214;
    reg node1215;
    reg node1216_r;
    reg node1216_l;
    reg node1217_r;
    reg node1217_l;
    reg node1218_r;
    reg node1218_l;
    reg node1219_r;
    reg node1219_l;
    reg node1220;
    reg node1221;
    reg node1222_r;
    reg node1222_l;
    reg node1223;
    reg node1224;
    reg node1225_r;
    reg node1225_l;
    reg node1226_r;
    reg node1226_l;
    reg node1227;
    reg node1228;
    reg node1229_r;
    reg node1229_l;
    reg node1230;
    reg node1231;
    reg node1232_r;
    reg node1232_l;
    reg node1233_r;
    reg node1233_l;
    reg node1234_r;
    reg node1234_l;
    reg node1235;
    reg node1236;
    reg node1237_r;
    reg node1237_l;
    reg node1238;
    reg node1239;
    reg node1240_r;
    reg node1240_l;
    reg node1241_r;
    reg node1241_l;
    reg node1242;
    reg node1243;
    reg node1244_r;
    reg node1244_l;
    reg node1245;
    reg node1246;
    reg node1247_r;
    reg node1247_l;
    reg node1248_r;
    reg node1248_l;
    reg node1249_r;
    reg node1249_l;
    reg node1250_r;
    reg node1250_l;
    reg node1251_r;
    reg node1251_l;
    reg node1252;
    reg node1253;
    reg node1254_r;
    reg node1254_l;
    reg node1255;
    reg node1256;
    reg node1257_r;
    reg node1257_l;
    reg node1258_r;
    reg node1258_l;
    reg node1259;
    reg node1260;
    reg node1261_r;
    reg node1261_l;
    reg node1262;
    reg node1263;
    reg node1264_r;
    reg node1264_l;
    reg node1265;
    reg node1266_r;
    reg node1266_l;
    reg node1267;
    reg node1268;
    reg node1269_r;
    reg node1269_l;
    reg node1270_r;
    reg node1270_l;
    reg node1271_r;
    reg node1271_l;
    reg node1272_r;
    reg node1272_l;
    reg node1273;
    reg node1274;
    reg node1275_r;
    reg node1275_l;
    reg node1276;
    reg node1277;
    reg node1278_r;
    reg node1278_l;
    reg node1279;
    reg node1280_r;
    reg node1280_l;
    reg node1281;
    reg node1282;
    reg node1283_r;
    reg node1283_l;
    reg node1284_r;
    reg node1284_l;
    reg node1285_r;
    reg node1285_l;
    reg node1286;
    reg node1287;
    reg node1288;
    reg node1289_r;
    reg node1289_l;
    reg node1290_r;
    reg node1290_l;
    reg node1291;
    reg node1292;
    reg node1293_r;
    reg node1293_l;
    reg node1294;
    reg node1295;
    reg node1296_r;
    reg node1296_l;
    reg node1297_r;
    reg node1297_l;
    reg node1298_r;
    reg node1298_l;
    reg node1299_r;
    reg node1299_l;
    reg node1300_r;
    reg node1300_l;
    reg node1301_r;
    reg node1301_l;
    reg node1302_r;
    reg node1302_l;
    reg node1303_r;
    reg node1303_l;
    reg node1304;
    reg node1305;
    reg node1306_r;
    reg node1306_l;
    reg node1307;
    reg node1308;
    reg node1309_r;
    reg node1309_l;
    reg node1310_r;
    reg node1310_l;
    reg node1311;
    reg node1312;
    reg node1313_r;
    reg node1313_l;
    reg node1314;
    reg node1315;
    reg node1316_r;
    reg node1316_l;
    reg node1317_r;
    reg node1317_l;
    reg node1318_r;
    reg node1318_l;
    reg node1319;
    reg node1320;
    reg node1321_r;
    reg node1321_l;
    reg node1322;
    reg node1323;
    reg node1324_r;
    reg node1324_l;
    reg node1325_r;
    reg node1325_l;
    reg node1326;
    reg node1327;
    reg node1328_r;
    reg node1328_l;
    reg node1329;
    reg node1330;
    reg node1331_r;
    reg node1331_l;
    reg node1332_r;
    reg node1332_l;
    reg node1333_r;
    reg node1333_l;
    reg node1334;
    reg node1335;
    reg node1336_r;
    reg node1336_l;
    reg node1337_r;
    reg node1337_l;
    reg node1338;
    reg node1339;
    reg node1340;
    reg node1341_r;
    reg node1341_l;
    reg node1342;
    reg node1343_r;
    reg node1343_l;
    reg node1344;
    reg node1345;
    reg node1346_r;
    reg node1346_l;
    reg node1347_r;
    reg node1347_l;
    reg node1348_r;
    reg node1348_l;
    reg node1349_r;
    reg node1349_l;
    reg node1350;
    reg node1351;
    reg node1352_r;
    reg node1352_l;
    reg node1353_r;
    reg node1353_l;
    reg node1354;
    reg node1355;
    reg node1356;
    reg node1357_r;
    reg node1357_l;
    reg node1358_r;
    reg node1358_l;
    reg node1359;
    reg node1360;
    reg node1361;
    reg node1362_r;
    reg node1362_l;
    reg node1363;
    reg node1364;
    reg node1365_r;
    reg node1365_l;
    reg node1366_r;
    reg node1366_l;
    reg node1367_r;
    reg node1367_l;
    reg node1368_r;
    reg node1368_l;
    reg node1369_r;
    reg node1369_l;
    reg node1370_r;
    reg node1370_l;
    reg node1371;
    reg node1372;
    reg node1373;
    reg node1374_r;
    reg node1374_l;
    reg node1375_r;
    reg node1375_l;
    reg node1376;
    reg node1377;
    reg node1378_r;
    reg node1378_l;
    reg node1379;
    reg node1380;
    reg node1381_r;
    reg node1381_l;
    reg node1382_r;
    reg node1382_l;
    reg node1383_r;
    reg node1383_l;
    reg node1384;
    reg node1385;
    reg node1386;
    reg node1387_r;
    reg node1387_l;
    reg node1388;
    reg node1389;
    reg node1390_r;
    reg node1390_l;
    reg node1391_r;
    reg node1391_l;
    reg node1392_r;
    reg node1392_l;
    reg node1393_r;
    reg node1393_l;
    reg node1394;
    reg node1395;
    reg node1396_r;
    reg node1396_l;
    reg node1397;
    reg node1398;
    reg node1399_r;
    reg node1399_l;
    reg node1400_r;
    reg node1400_l;
    reg node1401;
    reg node1402;
    reg node1403_r;
    reg node1403_l;
    reg node1404;
    reg node1405;
    reg node1406_r;
    reg node1406_l;
    reg node1407_r;
    reg node1407_l;
    reg node1408_r;
    reg node1408_l;
    reg node1409;
    reg node1410;
    reg node1411_r;
    reg node1411_l;
    reg node1412;
    reg node1413;
    reg node1414_r;
    reg node1414_l;
    reg node1415_r;
    reg node1415_l;
    reg node1416;
    reg node1417;
    reg node1418;
    reg node1419_r;
    reg node1419_l;
    reg node1420_r;
    reg node1420_l;
    reg node1421_r;
    reg node1421_l;
    reg node1422_r;
    reg node1422_l;
    reg node1423_r;
    reg node1423_l;
    reg node1424;
    reg node1425;
    reg node1426_r;
    reg node1426_l;
    reg node1427;
    reg node1428;
    reg node1429_r;
    reg node1429_l;
    reg node1430_r;
    reg node1430_l;
    reg node1431;
    reg node1432;
    reg node1433_r;
    reg node1433_l;
    reg node1434;
    reg node1435;
    reg node1436_r;
    reg node1436_l;
    reg node1437_r;
    reg node1437_l;
    reg node1438_r;
    reg node1438_l;
    reg node1439;
    reg node1440;
    reg node1441_r;
    reg node1441_l;
    reg node1442;
    reg node1443;
    reg node1444_r;
    reg node1444_l;
    reg node1445_r;
    reg node1445_l;
    reg node1446;
    reg node1447;
    reg node1448_r;
    reg node1448_l;
    reg node1449;
    reg node1450;
    reg node1451_r;
    reg node1451_l;
    reg node1452_r;
    reg node1452_l;
    reg node1453_r;
    reg node1453_l;
    reg node1454_r;
    reg node1454_l;
    reg node1455;
    reg node1456;
    reg node1457;
    reg node1458_r;
    reg node1458_l;
    reg node1459_r;
    reg node1459_l;
    reg node1460;
    reg node1461;
    reg node1462_r;
    reg node1462_l;
    reg node1463;
    reg node1464;
    reg node1465_r;
    reg node1465_l;
    reg node1466_r;
    reg node1466_l;
    reg node1467_r;
    reg node1467_l;
    reg node1468;
    reg node1469;
    reg node1470_r;
    reg node1470_l;
    reg node1471;
    reg node1472;
    reg node1473_r;
    reg node1473_l;
    reg node1474;
    reg node1475_r;
    reg node1475_l;
    reg node1476;
    reg node1477;
    reg node1478_r;
    reg node1478_l;
    reg node1479_r;
    reg node1479_l;
    reg node1480_r;
    reg node1480_l;
    reg node1481_r;
    reg node1481_l;
    reg node1482_r;
    reg node1482_l;
    reg node1483_r;
    reg node1483_l;
    reg node1484_r;
    reg node1484_l;
    reg node1485;
    reg node1486;
    reg node1487_r;
    reg node1487_l;
    reg node1488;
    reg node1489;
    reg node1490_r;
    reg node1490_l;
    reg node1491_r;
    reg node1491_l;
    reg node1492;
    reg node1493;
    reg node1494_r;
    reg node1494_l;
    reg node1495;
    reg node1496;
    reg node1497_r;
    reg node1497_l;
    reg node1498_r;
    reg node1498_l;
    reg node1499_r;
    reg node1499_l;
    reg node1500;
    reg node1501;
    reg node1502_r;
    reg node1502_l;
    reg node1503;
    reg node1504;
    reg node1505_r;
    reg node1505_l;
    reg node1506_r;
    reg node1506_l;
    reg node1507;
    reg node1508;
    reg node1509;
    reg node1510_r;
    reg node1510_l;
    reg node1511_r;
    reg node1511_l;
    reg node1512_r;
    reg node1512_l;
    reg node1513_r;
    reg node1513_l;
    reg node1514;
    reg node1515;
    reg node1516_r;
    reg node1516_l;
    reg node1517;
    reg node1518;
    reg node1519_r;
    reg node1519_l;
    reg node1520_r;
    reg node1520_l;
    reg node1521;
    reg node1522;
    reg node1523_r;
    reg node1523_l;
    reg node1524;
    reg node1525;
    reg node1526_r;
    reg node1526_l;
    reg node1527_r;
    reg node1527_l;
    reg node1528_r;
    reg node1528_l;
    reg node1529;
    reg node1530;
    reg node1531_r;
    reg node1531_l;
    reg node1532;
    reg node1533;
    reg node1534;
    reg node1535_r;
    reg node1535_l;
    reg node1536_r;
    reg node1536_l;
    reg node1537_r;
    reg node1537_l;
    reg node1538_r;
    reg node1538_l;
    reg node1539_r;
    reg node1539_l;
    reg node1540;
    reg node1541;
    reg node1542_r;
    reg node1542_l;
    reg node1543;
    reg node1544;
    reg node1545_r;
    reg node1545_l;
    reg node1546_r;
    reg node1546_l;
    reg node1547;
    reg node1548;
    reg node1549_r;
    reg node1549_l;
    reg node1550;
    reg node1551;
    reg node1552_r;
    reg node1552_l;
    reg node1553_r;
    reg node1553_l;
    reg node1554_r;
    reg node1554_l;
    reg node1555;
    reg node1556;
    reg node1557_r;
    reg node1557_l;
    reg node1558;
    reg node1559;
    reg node1560_r;
    reg node1560_l;
    reg node1561_r;
    reg node1561_l;
    reg node1562;
    reg node1563;
    reg node1564_r;
    reg node1564_l;
    reg node1565;
    reg node1566;
    reg node1567_r;
    reg node1567_l;
    reg node1568_r;
    reg node1568_l;
    reg node1569_r;
    reg node1569_l;
    reg node1570_r;
    reg node1570_l;
    reg node1571;
    reg node1572;
    reg node1573_r;
    reg node1573_l;
    reg node1574;
    reg node1575;
    reg node1576_r;
    reg node1576_l;
    reg node1577_r;
    reg node1577_l;
    reg node1578;
    reg node1579;
    reg node1580_r;
    reg node1580_l;
    reg node1581;
    reg node1582;
    reg node1583_r;
    reg node1583_l;
    reg node1584_r;
    reg node1584_l;
    reg node1585_r;
    reg node1585_l;
    reg node1586;
    reg node1587;
    reg node1588_r;
    reg node1588_l;
    reg node1589;
    reg node1590;
    reg node1591_r;
    reg node1591_l;
    reg node1592;
    reg node1593;
    reg node1594_r;
    reg node1594_l;
    reg node1595_r;
    reg node1595_l;
    reg node1596_r;
    reg node1596_l;
    reg node1597_r;
    reg node1597_l;
    reg node1598_r;
    reg node1598_l;
    reg node1599_r;
    reg node1599_l;
    reg node1600;
    reg node1601;
    reg node1602_r;
    reg node1602_l;
    reg node1603;
    reg node1604;
    reg node1605_r;
    reg node1605_l;
    reg node1606_r;
    reg node1606_l;
    reg node1607;
    reg node1608;
    reg node1609;
    reg node1610_r;
    reg node1610_l;
    reg node1611_r;
    reg node1611_l;
    reg node1612_r;
    reg node1612_l;
    reg node1613;
    reg node1614;
    reg node1615_r;
    reg node1615_l;
    reg node1616;
    reg node1617;
    reg node1618_r;
    reg node1618_l;
    reg node1619;
    reg node1620;
    reg node1621_r;
    reg node1621_l;
    reg node1622_r;
    reg node1622_l;
    reg node1623_r;
    reg node1623_l;
    reg node1624_r;
    reg node1624_l;
    reg node1625;
    reg node1626;
    reg node1627_r;
    reg node1627_l;
    reg node1628;
    reg node1629;
    reg node1630_r;
    reg node1630_l;
    reg node1631;
    reg node1632_r;
    reg node1632_l;
    reg node1633;
    reg node1634;
    reg node1635_r;
    reg node1635_l;
    reg node1636_r;
    reg node1636_l;
    reg node1637_r;
    reg node1637_l;
    reg node1638;
    reg node1639;
    reg node1640_r;
    reg node1640_l;
    reg node1641;
    reg node1642;
    reg node1643_r;
    reg node1643_l;
    reg node1644_r;
    reg node1644_l;
    reg node1645;
    reg node1646;
    reg node1647;
    reg node1648_r;
    reg node1648_l;
    reg node1649_r;
    reg node1649_l;
    reg node1650_r;
    reg node1650_l;
    reg node1651_r;
    reg node1651_l;
    reg node1652_r;
    reg node1652_l;
    reg node1653;
    reg node1654;
    reg node1655_r;
    reg node1655_l;
    reg node1656;
    reg node1657;
    reg node1658_r;
    reg node1658_l;
    reg node1659_r;
    reg node1659_l;
    reg node1660;
    reg node1661;
    reg node1662_r;
    reg node1662_l;
    reg node1663;
    reg node1664;
    reg node1665_r;
    reg node1665_l;
    reg node1666_r;
    reg node1666_l;
    reg node1667_r;
    reg node1667_l;
    reg node1668;
    reg node1669;
    reg node1670;
    reg node1671_r;
    reg node1671_l;
    reg node1672_r;
    reg node1672_l;
    reg node1673;
    reg node1674;
    reg node1675;
    reg node1676_r;
    reg node1676_l;
    reg node1677_r;
    reg node1677_l;
    reg node1678_r;
    reg node1678_l;
    reg node1679_r;
    reg node1679_l;
    reg node1680;
    reg node1681;
    reg node1682_r;
    reg node1682_l;
    reg node1683;
    reg node1684;
    reg node1685_r;
    reg node1685_l;
    reg node1686_r;
    reg node1686_l;
    reg node1687;
    reg node1688;
    reg node1689_r;
    reg node1689_l;
    reg node1690;
    reg node1691;
    reg node1692_r;
    reg node1692_l;
    reg node1693_r;
    reg node1693_l;
    reg node1694_r;
    reg node1694_l;
    reg node1695;
    reg node1696;
    reg node1697_r;
    reg node1697_l;
    reg node1698;
    reg node1699;
    reg node1700_r;
    reg node1700_l;
    reg node1701_r;
    reg node1701_l;
    reg node1702;
    reg node1703;
    reg node1704_r;
    reg node1704_l;
    reg node1705;
    reg node1706;
    reg result0;
    reg result1;
    reg result2;
    reg result3;
    reg result4;
    reg result5;
    reg result6;
    reg result7;
    reg result8;
    reg result9;

    begin
      node0_r = pixel[456];
      node0_l = ~pixel[456];
      node1_r = node0_l & pixel[290];
      node1_l = node0_l & ~pixel[290];
      node2_r = node1_l & pixel[488];
      node2_l = node1_l & ~pixel[488];
      node3_r = node2_l & pixel[655];
      node3_l = node2_l & ~pixel[655];
      node4_r = node3_l & pixel[598];
      node4_l = node3_l & ~pixel[598];
      node5_r = node4_l & pixel[438];
      node5_l = node4_l & ~pixel[438];
      node6_r = node5_l & pixel[353];
      node6_l = node5_l & ~pixel[353];
      node7_r = node6_l & pixel[490];
      node7_l = node6_l & ~pixel[490];
      node8_r = node7_l & pixel[373];
      node8_l = node7_l & ~pixel[373];
      node9_r = node8_l & pixel[712];
      node9_l = node8_l & ~pixel[712];
      node10 = node9_l;
      node11 = node9_r;
      node12_r = node8_r & pixel[104];
      node12_l = node8_r & ~pixel[104];
      node13 = node12_l;
      node14 = node12_r;
      node15_r = node7_r & pixel[406];
      node15_l = node7_r & ~pixel[406];
      node16_r = node15_l & pixel[433];
      node16_l = node15_l & ~pixel[433];
      node17 = node16_l;
      node18 = node16_r;
      node19_r = node15_r & pixel[325];
      node19_l = node15_r & ~pixel[325];
      node20 = node19_l;
      node21 = node19_r;
      node22_r = node6_r & pixel[454];
      node22_l = node6_r & ~pixel[454];
      node23_r = node22_l & pixel[344];
      node23_l = node22_l & ~pixel[344];
      node24_r = node23_l & pixel[203];
      node24_l = node23_l & ~pixel[203];
      node25 = node24_l;
      node26 = node24_r;
      node27_r = node23_r & pixel[551];
      node27_l = node23_r & ~pixel[551];
      node28 = node27_l;
      node29 = node27_r;
      node30_r = node22_r & pixel[400];
      node30_l = node22_r & ~pixel[400];
      node31_r = node30_l & pixel[468];
      node31_l = node30_l & ~pixel[468];
      node32 = node31_l;
      node33 = node31_r;
      node34_r = node30_r & pixel[184];
      node34_l = node30_r & ~pixel[184];
      node35 = node34_l;
      node36 = node34_r;
      node37_r = node5_r & pixel[235];
      node37_l = node5_r & ~pixel[235];
      node38_r = node37_l & pixel[181];
      node38_l = node37_l & ~pixel[181];
      node39_r = node38_l & pixel[540];
      node39_l = node38_l & ~pixel[540];
      node40_r = node39_l & pixel[102];
      node40_l = node39_l & ~pixel[102];
      node41 = node40_l;
      node42 = node40_r;
      node43_r = node39_r & pixel[368];
      node43_l = node39_r & ~pixel[368];
      node44 = node43_l;
      node45 = node43_r;
      node46_r = node38_r & pixel[491];
      node46_l = node38_r & ~pixel[491];
      node47_r = node46_l & pixel[342];
      node47_l = node46_l & ~pixel[342];
      node48 = node47_l;
      node49 = node47_r;
      node50_r = node46_r & pixel[260];
      node50_l = node46_r & ~pixel[260];
      node51 = node50_l;
      node52 = node50_r;
      node53_r = node37_r & pixel[607];
      node53_l = node37_r & ~pixel[607];
      node54_r = node53_l & pixel[432];
      node54_l = node53_l & ~pixel[432];
      node55_r = node54_l & pixel[375];
      node55_l = node54_l & ~pixel[375];
      node56 = node55_l;
      node57 = node55_r;
      node58_r = node54_r & pixel[688];
      node58_l = node54_r & ~pixel[688];
      node59 = node58_l;
      node60 = node58_r;
      node61_r = node53_r & pixel[322];
      node61_l = node53_r & ~pixel[322];
      node62_r = node61_l & pixel[601];
      node62_l = node61_l & ~pixel[601];
      node63 = node62_l;
      node64 = node62_r;
      node65_r = node61_r & pixel[720];
      node65_l = node61_r & ~pixel[720];
      node66 = node65_l;
      node67 = node65_r;
      node68_r = node4_r & pixel[220];
      node68_l = node4_r & ~pixel[220];
      node69_r = node68_l & pixel[292];
      node69_l = node68_l & ~pixel[292];
      node70_r = node69_l & pixel[359];
      node70_l = node69_l & ~pixel[359];
      node71_r = node70_l & pixel[522];
      node71_l = node70_l & ~pixel[522];
      node72_r = node71_l & pixel[514];
      node72_l = node71_l & ~pixel[514];
      node73 = node72_l;
      node74 = node72_r;
      node75_r = node71_r & pixel[379];
      node75_l = node71_r & ~pixel[379];
      node76 = node75_l;
      node77 = node75_r;
      node78_r = node70_r & pixel[463];
      node78_l = node70_r & ~pixel[463];
      node79_r = node78_l & pixel[405];
      node79_l = node78_l & ~pixel[405];
      node80 = node79_l;
      node81 = node79_r;
      node82_r = node78_r & pixel[161];
      node82_l = node78_r & ~pixel[161];
      node83 = node82_l;
      node84 = node82_r;
      node85_r = node69_r & pixel[247];
      node85_l = node69_r & ~pixel[247];
      node86_r = node85_l & pixel[538];
      node86_l = node85_l & ~pixel[538];
      node87_r = node86_l & pixel[568];
      node87_l = node86_l & ~pixel[568];
      node88 = node87_l;
      node89 = node87_r;
      node90_r = node86_r & pixel[535];
      node90_l = node86_r & ~pixel[535];
      node91 = node90_l;
      node92 = node90_r;
      node93_r = node85_r & pixel[270];
      node93_l = node85_r & ~pixel[270];
      node94_r = node93_l & pixel[237];
      node94_l = node93_l & ~pixel[237];
      node95 = node94_l;
      node96 = node94_r;
      node97_r = node93_r & pixel[432];
      node97_l = node93_r & ~pixel[432];
      node98 = node97_l;
      node99 = node97_r;
      node100_r = node68_r & pixel[355];
      node100_l = node68_r & ~pixel[355];
      node101_r = node100_l & pixel[426];
      node101_l = node100_l & ~pixel[426];
      node102 = node101_l;
      node103_r = node101_r & pixel[407];
      node103_l = node101_r & ~pixel[407];
      node104_r = node103_l & pixel[210];
      node104_l = node103_l & ~pixel[210];
      node105 = node104_l;
      node106 = node104_r;
      node107 = node103_r;
      node108_r = node100_r & pixel[211];
      node108_l = node100_r & ~pixel[211];
      node109 = node108_l;
      node110_r = node108_r & pixel[709];
      node110_l = node108_r & ~pixel[709];
      node111 = node110_l;
      node112 = node110_r;
      node113_r = node3_r & pixel[711];
      node113_l = node3_r & ~pixel[711];
      node114_r = node113_l & pixel[325];
      node114_l = node113_l & ~pixel[325];
      node115_r = node114_l & pixel[217];
      node115_l = node114_l & ~pixel[217];
      node116_r = node115_l & pixel[378];
      node116_l = node115_l & ~pixel[378];
      node117_r = node116_l & pixel[455];
      node117_l = node116_l & ~pixel[455];
      node118_r = node117_l & pixel[324];
      node118_l = node117_l & ~pixel[324];
      node119 = node118_l;
      node120 = node118_r;
      node121_r = node117_r & pixel[409];
      node121_l = node117_r & ~pixel[409];
      node122 = node121_l;
      node123 = node121_r;
      node124_r = node116_r & pixel[263];
      node124_l = node116_r & ~pixel[263];
      node125_r = node124_l & pixel[344];
      node125_l = node124_l & ~pixel[344];
      node126 = node125_l;
      node127 = node125_r;
      node128_r = node124_r & pixel[206];
      node128_l = node124_r & ~pixel[206];
      node129 = node128_l;
      node130 = node128_r;
      node131_r = node115_r & pixel[259];
      node131_l = node115_r & ~pixel[259];
      node132_r = node131_l & pixel[148];
      node132_l = node131_l & ~pixel[148];
      node133_r = node132_l & pixel[329];
      node133_l = node132_l & ~pixel[329];
      node134 = node133_l;
      node135 = node133_r;
      node136_r = node132_r & pixel[125];
      node136_l = node132_r & ~pixel[125];
      node137 = node136_l;
      node138 = node136_r;
      node139_r = node131_r & pixel[455];
      node139_l = node131_r & ~pixel[455];
      node140_r = node139_l & pixel[328];
      node140_l = node139_l & ~pixel[328];
      node141 = node140_l;
      node142 = node140_r;
      node143_r = node139_r & pixel[192];
      node143_l = node139_r & ~pixel[192];
      node144 = node143_l;
      node145 = node143_r;
      node146_r = node114_r & pixel[153];
      node146_l = node114_r & ~pixel[153];
      node147_r = node146_l & pixel[620];
      node147_l = node146_l & ~pixel[620];
      node148_r = node147_l & pixel[490];
      node148_l = node147_l & ~pixel[490];
      node149_r = node148_l & pixel[319];
      node149_l = node148_l & ~pixel[319];
      node150 = node149_l;
      node151 = node149_r;
      node152_r = node148_r & pixel[436];
      node152_l = node148_r & ~pixel[436];
      node153 = node152_l;
      node154 = node152_r;
      node155_r = node147_r & pixel[184];
      node155_l = node147_r & ~pixel[184];
      node156_r = node155_l & pixel[150];
      node156_l = node155_l & ~pixel[150];
      node157 = node156_l;
      node158 = node156_r;
      node159 = node155_r;
      node160_r = node146_r & pixel[315];
      node160_l = node146_r & ~pixel[315];
      node161_r = node160_l & pixel[623];
      node161_l = node160_l & ~pixel[623];
      node162_r = node161_l & pixel[375];
      node162_l = node161_l & ~pixel[375];
      node163 = node162_l;
      node164 = node162_r;
      node165_r = node161_r & pixel[611];
      node165_l = node161_r & ~pixel[611];
      node166 = node165_l;
      node167 = node165_r;
      node168_r = node160_r & pixel[427];
      node168_l = node160_r & ~pixel[427];
      node169_r = node168_l & pixel[321];
      node169_l = node168_l & ~pixel[321];
      node170 = node169_l;
      node171 = node169_r;
      node172_r = node168_r & pixel[270];
      node172_l = node168_r & ~pixel[270];
      node173 = node172_l;
      node174 = node172_r;
      node175_r = node113_r & pixel[346];
      node175_l = node113_r & ~pixel[346];
      node176_r = node175_l & pixel[519];
      node176_l = node175_l & ~pixel[519];
      node177_r = node176_l & pixel[180];
      node177_l = node176_l & ~pixel[180];
      node178_r = node177_l & pixel[234];
      node178_l = node177_l & ~pixel[234];
      node179_r = node178_l & pixel[268];
      node179_l = node178_l & ~pixel[268];
      node180 = node179_l;
      node181 = node179_r;
      node182_r = node178_r & pixel[551];
      node182_l = node178_r & ~pixel[551];
      node183 = node182_l;
      node184 = node182_r;
      node185_r = node177_r & pixel[192];
      node185_l = node177_r & ~pixel[192];
      node186_r = node185_l & pixel[350];
      node186_l = node185_l & ~pixel[350];
      node187 = node186_l;
      node188 = node186_r;
      node189 = node185_r;
      node190_r = node176_r & pixel[376];
      node190_l = node176_r & ~pixel[376];
      node191_r = node190_l & pixel[377];
      node191_l = node190_l & ~pixel[377];
      node192_r = node191_l & pixel[458];
      node192_l = node191_l & ~pixel[458];
      node193 = node192_l;
      node194 = node192_r;
      node195_r = node191_r & pixel[545];
      node195_l = node191_r & ~pixel[545];
      node196 = node195_l;
      node197 = node195_r;
      node198_r = node190_r & pixel[180];
      node198_l = node190_r & ~pixel[180];
      node199_r = node198_l & pixel[207];
      node199_l = node198_l & ~pixel[207];
      node200 = node199_l;
      node201 = node199_r;
      node202_r = node198_r & pixel[381];
      node202_l = node198_r & ~pixel[381];
      node203 = node202_l;
      node204 = node202_r;
      node205_r = node175_r & pixel[546];
      node205_l = node175_r & ~pixel[546];
      node206_r = node205_l & pixel[248];
      node206_l = node205_l & ~pixel[248];
      node207_r = node206_l & pixel[209];
      node207_l = node206_l & ~pixel[209];
      node208 = node207_l;
      node209_r = node207_r & pixel[596];
      node209_l = node207_r & ~pixel[596];
      node210 = node209_l;
      node211 = node209_r;
      node212 = node206_r;
      node213_r = node205_r & pixel[690];
      node213_l = node205_r & ~pixel[690];
      node214_r = node213_l & pixel[404];
      node214_l = node213_l & ~pixel[404];
      node215_r = node214_l & pixel[379];
      node215_l = node214_l & ~pixel[379];
      node216 = node215_l;
      node217 = node215_r;
      node218_r = node214_r & pixel[240];
      node218_l = node214_r & ~pixel[240];
      node219 = node218_l;
      node220 = node218_r;
      node221 = node213_r;
      node222_r = node2_r & pixel[606];
      node222_l = node2_r & ~pixel[606];
      node223_r = node222_l & pixel[206];
      node223_l = node222_l & ~pixel[206];
      node224_r = node223_l & pixel[402];
      node224_l = node223_l & ~pixel[402];
      node225_r = node224_l & pixel[327];
      node225_l = node224_l & ~pixel[327];
      node226_r = node225_l & pixel[323];
      node226_l = node225_l & ~pixel[323];
      node227_r = node226_l & pixel[241];
      node227_l = node226_l & ~pixel[241];
      node228_r = node227_l & pixel[186];
      node228_l = node227_l & ~pixel[186];
      node229 = node228_l;
      node230 = node228_r;
      node231_r = node227_r & pixel[404];
      node231_l = node227_r & ~pixel[404];
      node232 = node231_l;
      node233 = node231_r;
      node234_r = node226_r & pixel[464];
      node234_l = node226_r & ~pixel[464];
      node235_r = node234_l & pixel[523];
      node235_l = node234_l & ~pixel[523];
      node236 = node235_l;
      node237 = node235_r;
      node238_r = node234_r & pixel[568];
      node238_l = node234_r & ~pixel[568];
      node239 = node238_l;
      node240 = node238_r;
      node241_r = node225_r & pixel[520];
      node241_l = node225_r & ~pixel[520];
      node242_r = node241_l & pixel[292];
      node242_l = node241_l & ~pixel[292];
      node243_r = node242_l & pixel[632];
      node243_l = node242_l & ~pixel[632];
      node244 = node243_l;
      node245 = node243_r;
      node246_r = node242_r & pixel[597];
      node246_l = node242_r & ~pixel[597];
      node247 = node246_l;
      node248 = node246_r;
      node249_r = node241_r & pixel[379];
      node249_l = node241_r & ~pixel[379];
      node250_r = node249_l & pixel[655];
      node250_l = node249_l & ~pixel[655];
      node251 = node250_l;
      node252 = node250_r;
      node253_r = node249_r & pixel[265];
      node253_l = node249_r & ~pixel[265];
      node254 = node253_l;
      node255 = node253_r;
      node256_r = node224_r & pixel[521];
      node256_l = node224_r & ~pixel[521];
      node257_r = node256_l & pixel[463];
      node257_l = node256_l & ~pixel[463];
      node258_r = node257_l & pixel[578];
      node258_l = node257_l & ~pixel[578];
      node259_r = node258_l & pixel[513];
      node259_l = node258_l & ~pixel[513];
      node260 = node259_l;
      node261 = node259_r;
      node262 = node258_r;
      node263_r = node257_r & pixel[541];
      node263_l = node257_r & ~pixel[541];
      node264_r = node263_l & pixel[240];
      node264_l = node263_l & ~pixel[240];
      node265 = node264_l;
      node266 = node264_r;
      node267_r = node263_r & pixel[187];
      node267_l = node263_r & ~pixel[187];
      node268 = node267_l;
      node269 = node267_r;
      node270_r = node256_r & pixel[241];
      node270_l = node256_r & ~pixel[241];
      node271_r = node270_l & pixel[270];
      node271_l = node270_l & ~pixel[270];
      node272_r = node271_l & pixel[303];
      node272_l = node271_l & ~pixel[303];
      node273 = node272_l;
      node274 = node272_r;
      node275_r = node271_r & pixel[264];
      node275_l = node271_r & ~pixel[264];
      node276 = node275_l;
      node277 = node275_r;
      node278_r = node270_r & pixel[219];
      node278_l = node270_r & ~pixel[219];
      node279_r = node278_l & pixel[325];
      node279_l = node278_l & ~pixel[325];
      node280 = node279_l;
      node281 = node279_r;
      node282_r = node278_r & pixel[684];
      node282_l = node278_r & ~pixel[684];
      node283 = node282_l;
      node284 = node282_r;
      node285_r = node223_r & pixel[126];
      node285_l = node223_r & ~pixel[126];
      node286_r = node285_l & pixel[158];
      node286_l = node285_l & ~pixel[158];
      node287_r = node286_l & pixel[242];
      node287_l = node286_l & ~pixel[242];
      node288_r = node287_l & pixel[544];
      node288_l = node287_l & ~pixel[544];
      node289_r = node288_l & pixel[602];
      node289_l = node288_l & ~pixel[602];
      node290 = node289_l;
      node291 = node289_r;
      node292_r = node288_r & pixel[524];
      node292_l = node288_r & ~pixel[524];
      node293 = node292_l;
      node294 = node292_r;
      node295_r = node287_r & pixel[154];
      node295_l = node287_r & ~pixel[154];
      node296_r = node295_l & pixel[344];
      node296_l = node295_l & ~pixel[344];
      node297 = node296_l;
      node298 = node296_r;
      node299_r = node295_r & pixel[522];
      node299_l = node295_r & ~pixel[522];
      node300 = node299_l;
      node301 = node299_r;
      node302_r = node286_r & pixel[603];
      node302_l = node286_r & ~pixel[603];
      node303_r = node302_l & pixel[313];
      node303_l = node302_l & ~pixel[313];
      node304_r = node303_l & pixel[266];
      node304_l = node303_l & ~pixel[266];
      node305 = node304_l;
      node306 = node304_r;
      node307_r = node303_r & pixel[152];
      node307_l = node303_r & ~pixel[152];
      node308 = node307_l;
      node309 = node307_r;
      node310_r = node302_r & pixel[540];
      node310_l = node302_r & ~pixel[540];
      node311_r = node310_l & pixel[542];
      node311_l = node310_l & ~pixel[542];
      node312 = node311_l;
      node313 = node311_r;
      node314_r = node310_r & pixel[178];
      node314_l = node310_r & ~pixel[178];
      node315 = node314_l;
      node316 = node314_r;
      node317_r = node285_r & pixel[376];
      node317_l = node285_r & ~pixel[376];
      node318_r = node317_l & pixel[317];
      node318_l = node317_l & ~pixel[317];
      node319_r = node318_l & pixel[272];
      node319_l = node318_l & ~pixel[272];
      node320 = node319_l;
      node321_r = node319_r & pixel[351];
      node321_l = node319_r & ~pixel[351];
      node322 = node321_l;
      node323 = node321_r;
      node324_r = node318_r & pixel[627];
      node324_l = node318_r & ~pixel[627];
      node325 = node324_l;
      node326 = node324_r;
      node327_r = node317_r & pixel[554];
      node327_l = node317_r & ~pixel[554];
      node328_r = node327_l & pixel[326];
      node328_l = node327_l & ~pixel[326];
      node329_r = node328_l & pixel[414];
      node329_l = node328_l & ~pixel[414];
      node330 = node329_l;
      node331 = node329_r;
      node332_r = node328_r & pixel[497];
      node332_l = node328_r & ~pixel[497];
      node333 = node332_l;
      node334 = node332_r;
      node335 = node327_r;
      node336_r = node222_r & pixel[543];
      node336_l = node222_r & ~pixel[543];
      node337_r = node336_l & pixel[551];
      node337_l = node336_l & ~pixel[551];
      node338_r = node337_l & pixel[297];
      node338_l = node337_l & ~pixel[297];
      node339_r = node338_l & pixel[458];
      node339_l = node338_l & ~pixel[458];
      node340_r = node339_l & pixel[373];
      node340_l = node339_l & ~pixel[373];
      node341_r = node340_l & pixel[631];
      node341_l = node340_l & ~pixel[631];
      node342 = node341_l;
      node343 = node341_r;
      node344 = node340_r;
      node345_r = node339_r & pixel[299];
      node345_l = node339_r & ~pixel[299];
      node346_r = node345_l & pixel[513];
      node346_l = node345_l & ~pixel[513];
      node347 = node346_l;
      node348 = node346_r;
      node349_r = node345_r & pixel[258];
      node349_l = node345_r & ~pixel[258];
      node350 = node349_l;
      node351 = node349_r;
      node352_r = node338_r & pixel[542];
      node352_l = node338_r & ~pixel[542];
      node353_r = node352_l & pixel[654];
      node353_l = node352_l & ~pixel[654];
      node354_r = node353_l & pixel[465];
      node354_l = node353_l & ~pixel[465];
      node355 = node354_l;
      node356 = node354_r;
      node357_r = node353_r & pixel[345];
      node357_l = node353_r & ~pixel[345];
      node358 = node357_l;
      node359 = node357_r;
      node360_r = node352_r & pixel[444];
      node360_l = node352_r & ~pixel[444];
      node361_r = node360_l & pixel[550];
      node361_l = node360_l & ~pixel[550];
      node362 = node361_l;
      node363 = node361_r;
      node364 = node360_r;
      node365_r = node337_r & pixel[209];
      node365_l = node337_r & ~pixel[209];
      node366_r = node365_l & pixel[344];
      node366_l = node365_l & ~pixel[344];
      node367_r = node366_l & pixel[487];
      node367_l = node366_l & ~pixel[487];
      node368 = node367_l;
      node369_r = node367_r & pixel[271];
      node369_l = node367_r & ~pixel[271];
      node370 = node369_l;
      node371 = node369_r;
      node372_r = node366_r & pixel[459];
      node372_l = node366_r & ~pixel[459];
      node373_r = node372_l & pixel[661];
      node373_l = node372_l & ~pixel[661];
      node374 = node373_l;
      node375 = node373_r;
      node376_r = node372_r & pixel[327];
      node376_l = node372_r & ~pixel[327];
      node377 = node376_l;
      node378 = node376_r;
      node379_r = node365_r & pixel[150];
      node379_l = node365_r & ~pixel[150];
      node380_r = node379_l & pixel[317];
      node380_l = node379_l & ~pixel[317];
      node381_r = node380_l & pixel[378];
      node381_l = node380_l & ~pixel[378];
      node382 = node381_l;
      node383 = node381_r;
      node384_r = node380_r & pixel[428];
      node384_l = node380_r & ~pixel[428];
      node385 = node384_l;
      node386 = node384_r;
      node387_r = node379_r & pixel[523];
      node387_l = node379_r & ~pixel[523];
      node388_r = node387_l & pixel[188];
      node388_l = node387_l & ~pixel[188];
      node389 = node388_l;
      node390 = node388_r;
      node391_r = node387_r & pixel[605];
      node391_l = node387_r & ~pixel[605];
      node392 = node391_l;
      node393 = node391_r;
      node394_r = node336_r & pixel[403];
      node394_l = node336_r & ~pixel[403];
      node395_r = node394_l & pixel[397];
      node395_l = node394_l & ~pixel[397];
      node396_r = node395_l & pixel[541];
      node396_l = node395_l & ~pixel[541];
      node397_r = node396_l & pixel[439];
      node397_l = node396_l & ~pixel[439];
      node398_r = node397_l & pixel[203];
      node398_l = node397_l & ~pixel[203];
      node399 = node398_l;
      node400 = node398_r;
      node401_r = node397_r & pixel[375];
      node401_l = node397_r & ~pixel[375];
      node402 = node401_l;
      node403 = node401_r;
      node404_r = node396_r & pixel[292];
      node404_l = node396_r & ~pixel[292];
      node405_r = node404_l & pixel[298];
      node405_l = node404_l & ~pixel[298];
      node406 = node405_l;
      node407 = node405_r;
      node408_r = node404_r & pixel[659];
      node408_l = node404_r & ~pixel[659];
      node409 = node408_l;
      node410 = node408_r;
      node411_r = node395_r & pixel[609];
      node411_l = node395_r & ~pixel[609];
      node412 = node411_l;
      node413_r = node411_r & pixel[262];
      node413_l = node411_r & ~pixel[262];
      node414_r = node413_l & pixel[695];
      node414_l = node413_l & ~pixel[695];
      node415 = node414_l;
      node416 = node414_r;
      node417 = node413_r;
      node418_r = node394_r & pixel[123];
      node418_l = node394_r & ~pixel[123];
      node419_r = node418_l & pixel[319];
      node419_l = node418_l & ~pixel[319];
      node420_r = node419_l & pixel[686];
      node420_l = node419_l & ~pixel[686];
      node421_r = node420_l & pixel[633];
      node421_l = node420_l & ~pixel[633];
      node422 = node421_l;
      node423 = node421_r;
      node424_r = node420_r & pixel[343];
      node424_l = node420_r & ~pixel[343];
      node425 = node424_l;
      node426 = node424_r;
      node427_r = node419_r & pixel[297];
      node427_l = node419_r & ~pixel[297];
      node428_r = node427_l & pixel[265];
      node428_l = node427_l & ~pixel[265];
      node429 = node428_l;
      node430 = node428_r;
      node431_r = node427_r & pixel[324];
      node431_l = node427_r & ~pixel[324];
      node432 = node431_l;
      node433 = node431_r;
      node434_r = node418_r & pixel[659];
      node434_l = node418_r & ~pixel[659];
      node435_r = node434_l & pixel[440];
      node435_l = node434_l & ~pixel[440];
      node436_r = node435_l & pixel[358];
      node436_l = node435_l & ~pixel[358];
      node437 = node436_l;
      node438 = node436_r;
      node439_r = node435_r & pixel[428];
      node439_l = node435_r & ~pixel[428];
      node440 = node439_l;
      node441 = node439_r;
      node442_r = node434_r & pixel[468];
      node442_l = node434_r & ~pixel[468];
      node443_r = node442_l & pixel[374];
      node443_l = node442_l & ~pixel[374];
      node444 = node443_l;
      node445 = node443_r;
      node446_r = node442_r & pixel[598];
      node446_l = node442_r & ~pixel[598];
      node447 = node446_l;
      node448 = node446_r;
      node449_r = node1_r & pixel[406];
      node449_l = node1_r & ~pixel[406];
      node450_r = node449_l & pixel[437];
      node450_l = node449_l & ~pixel[437];
      node451_r = node450_l & pixel[386];
      node451_l = node450_l & ~pixel[386];
      node452_r = node451_l & pixel[190];
      node452_l = node451_l & ~pixel[190];
      node453_r = node452_l & pixel[444];
      node453_l = node452_l & ~pixel[444];
      node454_r = node453_l & pixel[625];
      node454_l = node453_l & ~pixel[625];
      node455_r = node454_l & pixel[260];
      node455_l = node454_l & ~pixel[260];
      node456_r = node455_l & pixel[490];
      node456_l = node455_l & ~pixel[490];
      node457 = node456_l;
      node458 = node456_r;
      node459_r = node455_r & pixel[327];
      node459_l = node455_r & ~pixel[327];
      node460 = node459_l;
      node461 = node459_r;
      node462_r = node454_r & pixel[350];
      node462_l = node454_r & ~pixel[350];
      node463_r = node462_l & pixel[370];
      node463_l = node462_l & ~pixel[370];
      node464 = node463_l;
      node465 = node463_r;
      node466_r = node462_r & pixel[121];
      node466_l = node462_r & ~pixel[121];
      node467 = node466_l;
      node468 = node466_r;
      node469_r = node453_r & pixel[454];
      node469_l = node453_r & ~pixel[454];
      node470_r = node469_l & pixel[68];
      node470_l = node469_l & ~pixel[68];
      node471 = node470_l;
      node472 = node470_r;
      node473 = node469_r;
      node474_r = node452_r & pixel[129];
      node474_l = node452_r & ~pixel[129];
      node475_r = node474_l & pixel[402];
      node475_l = node474_l & ~pixel[402];
      node476_r = node475_l & pixel[599];
      node476_l = node475_l & ~pixel[599];
      node477_r = node476_l & pixel[656];
      node477_l = node476_l & ~pixel[656];
      node478 = node477_l;
      node479 = node477_r;
      node480_r = node476_r & pixel[680];
      node480_l = node476_r & ~pixel[680];
      node481 = node480_l;
      node482 = node480_r;
      node483_r = node475_r & pixel[346];
      node483_l = node475_r & ~pixel[346];
      node484_r = node483_l & pixel[378];
      node484_l = node483_l & ~pixel[378];
      node485 = node484_l;
      node486 = node484_r;
      node487_r = node483_r & pixel[686];
      node487_l = node483_r & ~pixel[686];
      node488 = node487_l;
      node489 = node487_r;
      node490_r = node474_r & pixel[375];
      node490_l = node474_r & ~pixel[375];
      node491_r = node490_l & pixel[191];
      node491_l = node490_l & ~pixel[191];
      node492_r = node491_l & pixel[382];
      node492_l = node491_l & ~pixel[382];
      node493 = node492_l;
      node494 = node492_r;
      node495 = node491_r;
      node496 = node490_r;
      node497_r = node451_r & pixel[510];
      node497_l = node451_r & ~pixel[510];
      node498_r = node497_l & pixel[626];
      node498_l = node497_l & ~pixel[626];
      node499_r = node498_l & pixel[543];
      node499_l = node498_l & ~pixel[543];
      node500_r = node499_l & pixel[523];
      node500_l = node499_l & ~pixel[523];
      node501_r = node500_l & pixel[429];
      node501_l = node500_l & ~pixel[429];
      node502 = node501_l;
      node503 = node501_r;
      node504_r = node500_r & pixel[658];
      node504_l = node500_r & ~pixel[658];
      node505 = node504_l;
      node506 = node504_r;
      node507_r = node499_r & pixel[634];
      node507_l = node499_r & ~pixel[634];
      node508_r = node507_l & pixel[515];
      node508_l = node507_l & ~pixel[515];
      node509 = node508_l;
      node510 = node508_r;
      node511 = node507_r;
      node512_r = node498_r & pixel[425];
      node512_l = node498_r & ~pixel[425];
      node513_r = node512_l & pixel[354];
      node513_l = node512_l & ~pixel[354];
      node514_r = node513_l & pixel[610];
      node514_l = node513_l & ~pixel[610];
      node515 = node514_l;
      node516 = node514_r;
      node517_r = node513_r & pixel[200];
      node517_l = node513_r & ~pixel[200];
      node518 = node517_l;
      node519 = node517_r;
      node520_r = node512_r & pixel[576];
      node520_l = node512_r & ~pixel[576];
      node521_r = node520_l & pixel[604];
      node521_l = node520_l & ~pixel[604];
      node522 = node521_l;
      node523 = node521_r;
      node524 = node520_r;
      node525_r = node497_r & pixel[135];
      node525_l = node497_r & ~pixel[135];
      node526_r = node525_l & pixel[778];
      node526_l = node525_l & ~pixel[778];
      node527_r = node526_l & pixel[718];
      node527_l = node526_l & ~pixel[718];
      node528_r = node527_l & pixel[453];
      node528_l = node527_l & ~pixel[453];
      node529 = node528_l;
      node530 = node528_r;
      node531 = node527_r;
      node532 = node526_r;
      node533 = node525_r;
      node534_r = node450_r & pixel[402];
      node534_l = node450_r & ~pixel[402];
      node535_r = node534_l & pixel[569];
      node535_l = node534_l & ~pixel[569];
      node536_r = node535_l & pixel[151];
      node536_l = node535_l & ~pixel[151];
      node537_r = node536_l & pixel[190];
      node537_l = node536_l & ~pixel[190];
      node538_r = node537_l & pixel[460];
      node538_l = node537_l & ~pixel[460];
      node539_r = node538_l & pixel[267];
      node539_l = node538_l & ~pixel[267];
      node540 = node539_l;
      node541 = node539_r;
      node542_r = node538_r & pixel[231];
      node542_l = node538_r & ~pixel[231];
      node543 = node542_l;
      node544 = node542_r;
      node545_r = node537_r & pixel[518];
      node545_l = node537_r & ~pixel[518];
      node546 = node545_l;
      node547_r = node545_r & pixel[651];
      node547_l = node545_r & ~pixel[651];
      node548 = node547_l;
      node549 = node547_r;
      node550_r = node536_r & pixel[461];
      node550_l = node536_r & ~pixel[461];
      node551_r = node550_l & pixel[464];
      node551_l = node550_l & ~pixel[464];
      node552_r = node551_l & pixel[554];
      node552_l = node551_l & ~pixel[554];
      node553 = node552_l;
      node554 = node552_r;
      node555_r = node551_r & pixel[347];
      node555_l = node551_r & ~pixel[347];
      node556 = node555_l;
      node557 = node555_r;
      node558_r = node550_r & pixel[190];
      node558_l = node550_r & ~pixel[190];
      node559_r = node558_l & pixel[636];
      node559_l = node558_l & ~pixel[636];
      node560 = node559_l;
      node561 = node559_r;
      node562 = node558_r;
      node563_r = node535_r & pixel[435];
      node563_l = node535_r & ~pixel[435];
      node564_r = node563_l & pixel[490];
      node564_l = node563_l & ~pixel[490];
      node565_r = node564_l & pixel[235];
      node565_l = node564_l & ~pixel[235];
      node566_r = node565_l & pixel[627];
      node566_l = node565_l & ~pixel[627];
      node567 = node566_l;
      node568 = node566_r;
      node569_r = node565_r & pixel[432];
      node569_l = node565_r & ~pixel[432];
      node570 = node569_l;
      node571 = node569_r;
      node572_r = node564_r & pixel[206];
      node572_l = node564_r & ~pixel[206];
      node573_r = node572_l & pixel[595];
      node573_l = node572_l & ~pixel[595];
      node574 = node573_l;
      node575 = node573_r;
      node576_r = node572_r & pixel[453];
      node576_l = node572_r & ~pixel[453];
      node577 = node576_l;
      node578 = node576_r;
      node579_r = node563_r & pixel[180];
      node579_l = node563_r & ~pixel[180];
      node580_r = node579_l & pixel[566];
      node580_l = node579_l & ~pixel[566];
      node581_r = node580_l & pixel[544];
      node581_l = node580_l & ~pixel[544];
      node582 = node581_l;
      node583 = node581_r;
      node584_r = node580_r & pixel[657];
      node584_l = node580_r & ~pixel[657];
      node585 = node584_l;
      node586 = node584_r;
      node587_r = node579_r & pixel[99];
      node587_l = node579_r & ~pixel[99];
      node588_r = node587_l & pixel[481];
      node588_l = node587_l & ~pixel[481];
      node589 = node588_l;
      node590 = node588_r;
      node591_r = node587_r & pixel[371];
      node591_l = node587_r & ~pixel[371];
      node592 = node591_l;
      node593 = node591_r;
      node594_r = node534_r & pixel[98];
      node594_l = node534_r & ~pixel[98];
      node595_r = node594_l & pixel[597];
      node595_l = node594_l & ~pixel[597];
      node596_r = node595_l & pixel[266];
      node596_l = node595_l & ~pixel[266];
      node597_r = node596_l & pixel[97];
      node597_l = node596_l & ~pixel[97];
      node598_r = node597_l & pixel[431];
      node598_l = node597_l & ~pixel[431];
      node599 = node598_l;
      node600 = node598_r;
      node601 = node597_r;
      node602_r = node596_r & pixel[489];
      node602_l = node596_r & ~pixel[489];
      node603_r = node602_l & pixel[430];
      node603_l = node602_l & ~pixel[430];
      node604 = node603_l;
      node605 = node603_r;
      node606_r = node602_r & pixel[654];
      node606_l = node602_r & ~pixel[654];
      node607 = node606_l;
      node608 = node606_r;
      node609_r = node595_r & pixel[494];
      node609_l = node595_r & ~pixel[494];
      node610_r = node609_l & pixel[295];
      node610_l = node609_l & ~pixel[295];
      node611_r = node610_l & pixel[569];
      node611_l = node610_l & ~pixel[569];
      node612 = node611_l;
      node613 = node611_r;
      node614_r = node610_r & pixel[329];
      node614_l = node610_r & ~pixel[329];
      node615 = node614_l;
      node616 = node614_r;
      node617_r = node609_r & pixel[489];
      node617_l = node609_r & ~pixel[489];
      node618_r = node617_l & pixel[491];
      node618_l = node617_l & ~pixel[491];
      node619 = node618_l;
      node620 = node618_r;
      node621_r = node617_r & pixel[514];
      node621_l = node617_r & ~pixel[514];
      node622 = node621_l;
      node623 = node621_r;
      node624_r = node594_r & pixel[627];
      node624_l = node594_r & ~pixel[627];
      node625 = node624_l;
      node626_r = node624_r & pixel[374];
      node626_l = node624_r & ~pixel[374];
      node627 = node626_l;
      node628_r = node626_r & pixel[607];
      node628_l = node626_r & ~pixel[607];
      node629_r = node628_l & pixel[542];
      node629_l = node628_l & ~pixel[542];
      node630 = node629_l;
      node631 = node629_r;
      node632 = node628_r;
      node633_r = node449_r & pixel[186];
      node633_l = node449_r & ~pixel[186];
      node634_r = node633_l & pixel[402];
      node634_l = node633_l & ~pixel[402];
      node635_r = node634_l & pixel[151];
      node635_l = node634_l & ~pixel[151];
      node636_r = node635_l & pixel[156];
      node636_l = node635_l & ~pixel[156];
      node637_r = node636_l & pixel[297];
      node637_l = node636_l & ~pixel[297];
      node638_r = node637_l & pixel[212];
      node638_l = node637_l & ~pixel[212];
      node639_r = node638_l & pixel[459];
      node639_l = node638_l & ~pixel[459];
      node640 = node639_l;
      node641 = node639_r;
      node642_r = node638_r & pixel[569];
      node642_l = node638_r & ~pixel[569];
      node643 = node642_l;
      node644 = node642_r;
      node645_r = node637_r & pixel[374];
      node645_l = node637_r & ~pixel[374];
      node646_r = node645_l & pixel[555];
      node646_l = node645_l & ~pixel[555];
      node647 = node646_l;
      node648 = node646_r;
      node649_r = node645_r & pixel[348];
      node649_l = node645_r & ~pixel[348];
      node650 = node649_l;
      node651 = node649_r;
      node652_r = node636_r & pixel[459];
      node652_l = node636_r & ~pixel[459];
      node653_r = node652_l & pixel[327];
      node653_l = node652_l & ~pixel[327];
      node654_r = node653_l & pixel[295];
      node654_l = node653_l & ~pixel[295];
      node655 = node654_l;
      node656 = node654_r;
      node657_r = node653_r & pixel[376];
      node657_l = node653_r & ~pixel[376];
      node658 = node657_l;
      node659 = node657_r;
      node660_r = node652_r & pixel[414];
      node660_l = node652_r & ~pixel[414];
      node661_r = node660_l & pixel[455];
      node661_l = node660_l & ~pixel[455];
      node662 = node661_l;
      node663 = node661_r;
      node664_r = node660_r & pixel[656];
      node664_l = node660_r & ~pixel[656];
      node665 = node664_l;
      node666 = node664_r;
      node667_r = node635_r & pixel[347];
      node667_l = node635_r & ~pixel[347];
      node668_r = node667_l & pixel[545];
      node668_l = node667_l & ~pixel[545];
      node669_r = node668_l & pixel[297];
      node669_l = node668_l & ~pixel[297];
      node670_r = node669_l & pixel[323];
      node670_l = node669_l & ~pixel[323];
      node671 = node670_l;
      node672 = node670_r;
      node673_r = node669_r & pixel[288];
      node673_l = node669_r & ~pixel[288];
      node674 = node673_l;
      node675 = node673_r;
      node676_r = node668_r & pixel[510];
      node676_l = node668_r & ~pixel[510];
      node677_r = node676_l & pixel[434];
      node677_l = node676_l & ~pixel[434];
      node678 = node677_l;
      node679 = node677_r;
      node680 = node676_r;
      node681_r = node667_r & pixel[460];
      node681_l = node667_r & ~pixel[460];
      node682_r = node681_l & pixel[491];
      node682_l = node681_l & ~pixel[491];
      node683_r = node682_l & pixel[321];
      node683_l = node682_l & ~pixel[321];
      node684 = node683_l;
      node685 = node683_r;
      node686_r = node682_r & pixel[241];
      node686_l = node682_r & ~pixel[241];
      node687 = node686_l;
      node688 = node686_r;
      node689_r = node681_r & pixel[575];
      node689_l = node681_r & ~pixel[575];
      node690_r = node689_l & pixel[633];
      node690_l = node689_l & ~pixel[633];
      node691 = node690_l;
      node692 = node690_r;
      node693_r = node689_r & pixel[486];
      node693_l = node689_r & ~pixel[486];
      node694 = node693_l;
      node695 = node693_r;
      node696_r = node634_r & pixel[567];
      node696_l = node634_r & ~pixel[567];
      node697_r = node696_l & pixel[241];
      node697_l = node696_l & ~pixel[241];
      node698_r = node697_l & pixel[271];
      node698_l = node697_l & ~pixel[271];
      node699_r = node698_l & pixel[459];
      node699_l = node698_l & ~pixel[459];
      node700_r = node699_l & pixel[352];
      node700_l = node699_l & ~pixel[352];
      node701 = node700_l;
      node702 = node700_r;
      node703_r = node699_r & pixel[660];
      node703_l = node699_r & ~pixel[660];
      node704 = node703_l;
      node705 = node703_r;
      node706_r = node698_r & pixel[383];
      node706_l = node698_r & ~pixel[383];
      node707_r = node706_l & pixel[605];
      node707_l = node706_l & ~pixel[605];
      node708 = node707_l;
      node709 = node707_r;
      node710_r = node706_r & pixel[148];
      node710_l = node706_r & ~pixel[148];
      node711 = node710_l;
      node712 = node710_r;
      node713_r = node697_r & pixel[516];
      node713_l = node697_r & ~pixel[516];
      node714_r = node713_l & pixel[409];
      node714_l = node713_l & ~pixel[409];
      node715_r = node714_l & pixel[628];
      node715_l = node714_l & ~pixel[628];
      node716 = node715_l;
      node717 = node715_r;
      node718_r = node714_r & pixel[154];
      node718_l = node714_r & ~pixel[154];
      node719 = node718_l;
      node720 = node718_r;
      node721_r = node713_r & pixel[635];
      node721_l = node713_r & ~pixel[635];
      node722_r = node721_l & pixel[240];
      node722_l = node721_l & ~pixel[240];
      node723 = node722_l;
      node724 = node722_r;
      node725_r = node721_r & pixel[543];
      node725_l = node721_r & ~pixel[543];
      node726 = node725_l;
      node727 = node725_r;
      node728_r = node696_r & pixel[180];
      node728_l = node696_r & ~pixel[180];
      node729_r = node728_l & pixel[487];
      node729_l = node728_l & ~pixel[487];
      node730_r = node729_l & pixel[460];
      node730_l = node729_l & ~pixel[460];
      node731_r = node730_l & pixel[206];
      node731_l = node730_l & ~pixel[206];
      node732 = node731_l;
      node733 = node731_r;
      node734_r = node730_r & pixel[381];
      node734_l = node730_r & ~pixel[381];
      node735 = node734_l;
      node736 = node734_r;
      node737_r = node729_r & pixel[486];
      node737_l = node729_r & ~pixel[486];
      node738 = node737_l;
      node739_r = node737_r & pixel[628];
      node739_l = node737_r & ~pixel[628];
      node740 = node739_l;
      node741 = node739_r;
      node742_r = node728_r & pixel[306];
      node742_l = node728_r & ~pixel[306];
      node743_r = node742_l & pixel[460];
      node743_l = node742_l & ~pixel[460];
      node744_r = node743_l & pixel[216];
      node744_l = node743_l & ~pixel[216];
      node745 = node744_l;
      node746 = node744_r;
      node747_r = node743_r & pixel[488];
      node747_l = node743_r & ~pixel[488];
      node748 = node747_l;
      node749 = node747_r;
      node750 = node742_r;
      node751_r = node633_r & pixel[271];
      node751_l = node633_r & ~pixel[271];
      node752_r = node751_l & pixel[518];
      node752_l = node751_l & ~pixel[518];
      node753_r = node752_l & pixel[653];
      node753_l = node752_l & ~pixel[653];
      node754_r = node753_l & pixel[160];
      node754_l = node753_l & ~pixel[160];
      node755_r = node754_l & pixel[656];
      node755_l = node754_l & ~pixel[656];
      node756_r = node755_l & pixel[211];
      node756_l = node755_l & ~pixel[211];
      node757 = node756_l;
      node758 = node756_r;
      node759_r = node755_r & pixel[543];
      node759_l = node755_r & ~pixel[543];
      node760 = node759_l;
      node761 = node759_r;
      node762_r = node754_r & pixel[296];
      node762_l = node754_r & ~pixel[296];
      node763_r = node762_l & pixel[487];
      node763_l = node762_l & ~pixel[487];
      node764 = node763_l;
      node765 = node763_r;
      node766_r = node762_r & pixel[575];
      node766_l = node762_r & ~pixel[575];
      node767 = node766_l;
      node768 = node766_r;
      node769_r = node753_r & pixel[246];
      node769_l = node753_r & ~pixel[246];
      node770_r = node769_l & pixel[122];
      node770_l = node769_l & ~pixel[122];
      node771_r = node770_l & pixel[300];
      node771_l = node770_l & ~pixel[300];
      node772 = node771_l;
      node773 = node771_r;
      node774_r = node770_r & pixel[158];
      node774_l = node770_r & ~pixel[158];
      node775 = node774_l;
      node776 = node774_r;
      node777_r = node769_r & pixel[302];
      node777_l = node769_r & ~pixel[302];
      node778_r = node777_l & pixel[328];
      node778_l = node777_l & ~pixel[328];
      node779 = node778_l;
      node780 = node778_r;
      node781_r = node777_r & pixel[489];
      node781_l = node777_r & ~pixel[489];
      node782 = node781_l;
      node783 = node781_r;
      node784_r = node752_r & pixel[162];
      node784_l = node752_r & ~pixel[162];
      node785_r = node784_l & pixel[272];
      node785_l = node784_l & ~pixel[272];
      node786_r = node785_l & pixel[543];
      node786_l = node785_l & ~pixel[543];
      node787_r = node786_l & pixel[381];
      node787_l = node786_l & ~pixel[381];
      node788 = node787_l;
      node789 = node787_r;
      node790_r = node786_r & pixel[684];
      node790_l = node786_r & ~pixel[684];
      node791 = node790_l;
      node792 = node790_r;
      node793_r = node785_r & pixel[572];
      node793_l = node785_r & ~pixel[572];
      node794_r = node793_l & pixel[427];
      node794_l = node793_l & ~pixel[427];
      node795 = node794_l;
      node796 = node794_r;
      node797_r = node793_r & pixel[659];
      node797_l = node793_r & ~pixel[659];
      node798 = node797_l;
      node799 = node797_r;
      node800_r = node784_r & pixel[486];
      node800_l = node784_r & ~pixel[486];
      node801_r = node800_l & pixel[480];
      node801_l = node800_l & ~pixel[480];
      node802_r = node801_l & pixel[204];
      node802_l = node801_l & ~pixel[204];
      node803 = node802_l;
      node804 = node802_r;
      node805_r = node801_r & pixel[516];
      node805_l = node801_r & ~pixel[516];
      node806 = node805_l;
      node807 = node805_r;
      node808_r = node800_r & pixel[460];
      node808_l = node800_r & ~pixel[460];
      node809 = node808_l;
      node810_r = node808_r & pixel[482];
      node810_l = node808_r & ~pixel[482];
      node811 = node810_l;
      node812 = node810_r;
      node813_r = node751_r & pixel[238];
      node813_l = node751_r & ~pixel[238];
      node814_r = node813_l & pixel[401];
      node814_l = node813_l & ~pixel[401];
      node815_r = node814_l & pixel[318];
      node815_l = node814_l & ~pixel[318];
      node816_r = node815_l & pixel[349];
      node816_l = node815_l & ~pixel[349];
      node817_r = node816_l & pixel[684];
      node817_l = node816_l & ~pixel[684];
      node818 = node817_l;
      node819 = node817_r;
      node820_r = node816_r & pixel[496];
      node820_l = node816_r & ~pixel[496];
      node821 = node820_l;
      node822 = node820_r;
      node823_r = node815_r & pixel[487];
      node823_l = node815_r & ~pixel[487];
      node824_r = node823_l & pixel[595];
      node824_l = node823_l & ~pixel[595];
      node825 = node824_l;
      node826 = node824_r;
      node827_r = node823_r & pixel[376];
      node827_l = node823_r & ~pixel[376];
      node828 = node827_l;
      node829 = node827_r;
      node830_r = node814_r & pixel[569];
      node830_l = node814_r & ~pixel[569];
      node831_r = node830_l & pixel[185];
      node831_l = node830_l & ~pixel[185];
      node832_r = node831_l & pixel[154];
      node832_l = node831_l & ~pixel[154];
      node833 = node832_l;
      node834 = node832_r;
      node835_r = node831_r & pixel[354];
      node835_l = node831_r & ~pixel[354];
      node836 = node835_l;
      node837 = node835_r;
      node838_r = node830_r & pixel[326];
      node838_l = node830_r & ~pixel[326];
      node839_r = node838_l & pixel[320];
      node839_l = node838_l & ~pixel[320];
      node840 = node839_l;
      node841 = node839_r;
      node842_r = node838_r & pixel[594];
      node842_l = node838_r & ~pixel[594];
      node843 = node842_l;
      node844 = node842_r;
      node845_r = node813_r & pixel[155];
      node845_l = node813_r & ~pixel[155];
      node846_r = node845_l & pixel[568];
      node846_l = node845_l & ~pixel[568];
      node847_r = node846_l & pixel[345];
      node847_l = node846_l & ~pixel[345];
      node848_r = node847_l & pixel[261];
      node848_l = node847_l & ~pixel[261];
      node849 = node848_l;
      node850 = node848_r;
      node851_r = node847_r & pixel[576];
      node851_l = node847_r & ~pixel[576];
      node852 = node851_l;
      node853 = node851_r;
      node854_r = node846_r & pixel[352];
      node854_l = node846_r & ~pixel[352];
      node855_r = node854_l & pixel[382];
      node855_l = node854_l & ~pixel[382];
      node856 = node855_l;
      node857 = node855_r;
      node858_r = node854_r & pixel[463];
      node858_l = node854_r & ~pixel[463];
      node859 = node858_l;
      node860 = node858_r;
      node861_r = node845_r & pixel[537];
      node861_l = node845_r & ~pixel[537];
      node862_r = node861_l & pixel[552];
      node862_l = node861_l & ~pixel[552];
      node863_r = node862_l & pixel[488];
      node863_l = node862_l & ~pixel[488];
      node864 = node863_l;
      node865 = node863_r;
      node866_r = node862_r & pixel[346];
      node866_l = node862_r & ~pixel[346];
      node867 = node866_l;
      node868 = node866_r;
      node869_r = node861_r & pixel[344];
      node869_l = node861_r & ~pixel[344];
      node870_r = node869_l & pixel[515];
      node870_l = node869_l & ~pixel[515];
      node871 = node870_l;
      node872 = node870_r;
      node873_r = node869_r & pixel[356];
      node873_l = node869_r & ~pixel[356];
      node874 = node873_l;
      node875 = node873_r;
      node876_r = node0_r & pixel[380];
      node876_l = node0_r & ~pixel[380];
      node877_r = node876_l & pixel[185];
      node877_l = node876_l & ~pixel[185];
      node878_r = node877_l & pixel[213];
      node878_l = node877_l & ~pixel[213];
      node879_r = node878_l & pixel[497];
      node879_l = node878_l & ~pixel[497];
      node880_r = node879_l & pixel[101];
      node880_l = node879_l & ~pixel[101];
      node881_r = node880_l & pixel[269];
      node881_l = node880_l & ~pixel[269];
      node882_r = node881_l & pixel[296];
      node882_l = node881_l & ~pixel[296];
      node883_r = node882_l & pixel[355];
      node883_l = node882_l & ~pixel[355];
      node884_r = node883_l & pixel[571];
      node884_l = node883_l & ~pixel[571];
      node885 = node884_l;
      node886 = node884_r;
      node887_r = node883_r & pixel[650];
      node887_l = node883_r & ~pixel[650];
      node888 = node887_l;
      node889 = node887_r;
      node890_r = node882_r & pixel[386];
      node890_l = node882_r & ~pixel[386];
      node891_r = node890_l & pixel[383];
      node891_l = node890_l & ~pixel[383];
      node892 = node891_l;
      node893 = node891_r;
      node894_r = node890_r & pixel[571];
      node894_l = node890_r & ~pixel[571];
      node895 = node894_l;
      node896 = node894_r;
      node897_r = node881_r & pixel[355];
      node897_l = node881_r & ~pixel[355];
      node898_r = node897_l & pixel[414];
      node898_l = node897_l & ~pixel[414];
      node899_r = node898_l & pixel[714];
      node899_l = node898_l & ~pixel[714];
      node900 = node899_l;
      node901 = node899_r;
      node902_r = node898_r & pixel[440];
      node902_l = node898_r & ~pixel[440];
      node903 = node902_l;
      node904 = node902_r;
      node905_r = node897_r & pixel[461];
      node905_l = node897_r & ~pixel[461];
      node906_r = node905_l & pixel[543];
      node906_l = node905_l & ~pixel[543];
      node907 = node906_l;
      node908 = node906_r;
      node909_r = node905_r & pixel[215];
      node909_l = node905_r & ~pixel[215];
      node910 = node909_l;
      node911 = node909_r;
      node912_r = node880_r & pixel[188];
      node912_l = node880_r & ~pixel[188];
      node913_r = node912_l & pixel[467];
      node913_l = node912_l & ~pixel[467];
      node914_r = node913_l & pixel[485];
      node914_l = node913_l & ~pixel[485];
      node915_r = node914_l & pixel[602];
      node915_l = node914_l & ~pixel[602];
      node916 = node915_l;
      node917 = node915_r;
      node918_r = node914_r & pixel[289];
      node918_l = node914_r & ~pixel[289];
      node919 = node918_l;
      node920 = node918_r;
      node921_r = node913_r & pixel[329];
      node921_l = node913_r & ~pixel[329];
      node922_r = node921_l & pixel[512];
      node922_l = node921_l & ~pixel[512];
      node923 = node922_l;
      node924 = node922_r;
      node925_r = node921_r & pixel[346];
      node925_l = node921_r & ~pixel[346];
      node926 = node925_l;
      node927 = node925_r;
      node928_r = node912_r & pixel[482];
      node928_l = node912_r & ~pixel[482];
      node929_r = node928_l & pixel[210];
      node929_l = node928_l & ~pixel[210];
      node930 = node929_l;
      node931_r = node929_r & pixel[405];
      node931_l = node929_r & ~pixel[405];
      node932 = node931_l;
      node933 = node931_r;
      node934_r = node928_r & pixel[293];
      node934_l = node928_r & ~pixel[293];
      node935_r = node934_l & pixel[415];
      node935_l = node934_l & ~pixel[415];
      node936 = node935_l;
      node937 = node935_r;
      node938_r = node934_r & pixel[322];
      node938_l = node934_r & ~pixel[322];
      node939 = node938_l;
      node940 = node938_r;
      node941_r = node879_r & pixel[272];
      node941_l = node879_r & ~pixel[272];
      node942_r = node941_l & pixel[409];
      node942_l = node941_l & ~pixel[409];
      node943_r = node942_l & pixel[577];
      node943_l = node942_l & ~pixel[577];
      node944_r = node943_l & pixel[345];
      node944_l = node943_l & ~pixel[345];
      node945_r = node944_l & pixel[684];
      node945_l = node944_l & ~pixel[684];
      node946 = node945_l;
      node947 = node945_r;
      node948_r = node944_r & pixel[512];
      node948_l = node944_r & ~pixel[512];
      node949 = node948_l;
      node950 = node948_r;
      node951_r = node943_r & pixel[100];
      node951_l = node943_r & ~pixel[100];
      node952_r = node951_l & pixel[432];
      node952_l = node951_l & ~pixel[432];
      node953 = node952_l;
      node954 = node952_r;
      node955_r = node951_r & pixel[549];
      node955_l = node951_r & ~pixel[549];
      node956 = node955_l;
      node957 = node955_r;
      node958_r = node942_r & pixel[324];
      node958_l = node942_r & ~pixel[324];
      node959_r = node958_l & pixel[270];
      node959_l = node958_l & ~pixel[270];
      node960_r = node959_l & pixel[275];
      node960_l = node959_l & ~pixel[275];
      node961 = node960_l;
      node962 = node960_r;
      node963_r = node959_r & pixel[499];
      node963_l = node959_r & ~pixel[499];
      node964 = node963_l;
      node965 = node963_r;
      node966_r = node958_r & pixel[183];
      node966_l = node958_r & ~pixel[183];
      node967_r = node966_l & pixel[437];
      node967_l = node966_l & ~pixel[437];
      node968 = node967_l;
      node969 = node967_r;
      node970_r = node966_r & pixel[379];
      node970_l = node966_r & ~pixel[379];
      node971 = node970_l;
      node972 = node970_r;
      node973_r = node941_r & pixel[359];
      node973_l = node941_r & ~pixel[359];
      node974_r = node973_l & pixel[269];
      node974_l = node973_l & ~pixel[269];
      node975_r = node974_l & pixel[129];
      node975_l = node974_l & ~pixel[129];
      node976_r = node975_l & pixel[92];
      node976_l = node975_l & ~pixel[92];
      node977 = node976_l;
      node978 = node976_r;
      node979_r = node975_r & pixel[438];
      node979_l = node975_r & ~pixel[438];
      node980 = node979_l;
      node981 = node979_r;
      node982_r = node974_r & pixel[178];
      node982_l = node974_r & ~pixel[178];
      node983_r = node982_l & pixel[543];
      node983_l = node982_l & ~pixel[543];
      node984 = node983_l;
      node985 = node983_r;
      node986_r = node982_r & pixel[659];
      node986_l = node982_r & ~pixel[659];
      node987 = node986_l;
      node988 = node986_r;
      node989_r = node973_r & pixel[93];
      node989_l = node973_r & ~pixel[93];
      node990_r = node989_l & pixel[639];
      node990_l = node989_l & ~pixel[639];
      node991_r = node990_l & pixel[454];
      node991_l = node990_l & ~pixel[454];
      node992 = node991_l;
      node993 = node991_r;
      node994 = node990_r;
      node995_r = node989_r & pixel[119];
      node995_l = node989_r & ~pixel[119];
      node996 = node995_l;
      node997_r = node995_r & pixel[348];
      node997_l = node995_r & ~pixel[348];
      node998 = node997_l;
      node999 = node997_r;
      node1000_r = node878_r & pixel[386];
      node1000_l = node878_r & ~pixel[386];
      node1001_r = node1000_l & pixel[626];
      node1001_l = node1000_l & ~pixel[626];
      node1002_r = node1001_l & pixel[218];
      node1002_l = node1001_l & ~pixel[218];
      node1003_r = node1002_l & pixel[686];
      node1003_l = node1002_l & ~pixel[686];
      node1004_r = node1003_l & pixel[554];
      node1004_l = node1003_l & ~pixel[554];
      node1005_r = node1004_l & pixel[539];
      node1005_l = node1004_l & ~pixel[539];
      node1006 = node1005_l;
      node1007 = node1005_r;
      node1008_r = node1004_r & pixel[341];
      node1008_l = node1004_r & ~pixel[341];
      node1009 = node1008_l;
      node1010 = node1008_r;
      node1011_r = node1003_r & pixel[460];
      node1011_l = node1003_r & ~pixel[460];
      node1012_r = node1011_l & pixel[344];
      node1012_l = node1011_l & ~pixel[344];
      node1013 = node1012_l;
      node1014 = node1012_r;
      node1015_r = node1011_r & pixel[465];
      node1015_l = node1011_r & ~pixel[465];
      node1016 = node1015_l;
      node1017 = node1015_r;
      node1018_r = node1002_r & pixel[632];
      node1018_l = node1002_r & ~pixel[632];
      node1019_r = node1018_l & pixel[565];
      node1019_l = node1018_l & ~pixel[565];
      node1020_r = node1019_l & pixel[467];
      node1020_l = node1019_l & ~pixel[467];
      node1021 = node1020_l;
      node1022 = node1020_r;
      node1023_r = node1019_r & pixel[409];
      node1023_l = node1019_r & ~pixel[409];
      node1024 = node1023_l;
      node1025 = node1023_r;
      node1026_r = node1018_r & pixel[313];
      node1026_l = node1018_r & ~pixel[313];
      node1027 = node1026_l;
      node1028 = node1026_r;
      node1029_r = node1001_r & pixel[385];
      node1029_l = node1001_r & ~pixel[385];
      node1030_r = node1029_l & pixel[154];
      node1030_l = node1029_l & ~pixel[154];
      node1031_r = node1030_l & pixel[248];
      node1031_l = node1030_l & ~pixel[248];
      node1032_r = node1031_l & pixel[658];
      node1032_l = node1031_l & ~pixel[658];
      node1033 = node1032_l;
      node1034 = node1032_r;
      node1035_r = node1031_r & pixel[438];
      node1035_l = node1031_r & ~pixel[438];
      node1036 = node1035_l;
      node1037 = node1035_r;
      node1038_r = node1030_r & pixel[193];
      node1038_l = node1030_r & ~pixel[193];
      node1039_r = node1038_l & pixel[518];
      node1039_l = node1038_l & ~pixel[518];
      node1040 = node1039_l;
      node1041 = node1039_r;
      node1042 = node1038_r;
      node1043_r = node1029_r & pixel[709];
      node1043_l = node1029_r & ~pixel[709];
      node1044_r = node1043_l & pixel[401];
      node1044_l = node1043_l & ~pixel[401];
      node1045_r = node1044_l & pixel[430];
      node1045_l = node1044_l & ~pixel[430];
      node1046 = node1045_l;
      node1047 = node1045_r;
      node1048_r = node1044_r & pixel[459];
      node1048_l = node1044_r & ~pixel[459];
      node1049 = node1048_l;
      node1050 = node1048_r;
      node1051_r = node1043_r & pixel[316];
      node1051_l = node1043_r & ~pixel[316];
      node1052 = node1051_l;
      node1053 = node1051_r;
      node1054_r = node1000_r & pixel[573];
      node1054_l = node1000_r & ~pixel[573];
      node1055_r = node1054_l & pixel[435];
      node1055_l = node1054_l & ~pixel[435];
      node1056_r = node1055_l & pixel[541];
      node1056_l = node1055_l & ~pixel[541];
      node1057_r = node1056_l & pixel[595];
      node1057_l = node1056_l & ~pixel[595];
      node1058_r = node1057_l & pixel[266];
      node1058_l = node1057_l & ~pixel[266];
      node1059 = node1058_l;
      node1060 = node1058_r;
      node1061 = node1057_r;
      node1062 = node1056_r;
      node1063_r = node1055_r & pixel[302];
      node1063_l = node1055_r & ~pixel[302];
      node1064_r = node1063_l & pixel[370];
      node1064_l = node1063_l & ~pixel[370];
      node1065 = node1064_l;
      node1066_r = node1064_r & pixel[653];
      node1066_l = node1064_r & ~pixel[653];
      node1067 = node1066_l;
      node1068 = node1066_r;
      node1069_r = node1063_r & pixel[186];
      node1069_l = node1063_r & ~pixel[186];
      node1070_r = node1069_l & pixel[494];
      node1070_l = node1069_l & ~pixel[494];
      node1071 = node1070_l;
      node1072 = node1070_r;
      node1073 = node1069_r;
      node1074_r = node1054_r & pixel[462];
      node1074_l = node1054_r & ~pixel[462];
      node1075_r = node1074_l & pixel[740];
      node1075_l = node1074_l & ~pixel[740];
      node1076_r = node1075_l & pixel[368];
      node1076_l = node1075_l & ~pixel[368];
      node1077_r = node1076_l & pixel[745];
      node1077_l = node1076_l & ~pixel[745];
      node1078 = node1077_l;
      node1079 = node1077_r;
      node1080_r = node1076_r & pixel[291];
      node1080_l = node1076_r & ~pixel[291];
      node1081 = node1080_l;
      node1082 = node1080_r;
      node1083 = node1075_r;
      node1084_r = node1074_r & pixel[708];
      node1084_l = node1074_r & ~pixel[708];
      node1085_r = node1084_l & pixel[176];
      node1085_l = node1084_l & ~pixel[176];
      node1086_r = node1085_l & pixel[626];
      node1086_l = node1085_l & ~pixel[626];
      node1087 = node1086_l;
      node1088 = node1086_r;
      node1089 = node1085_r;
      node1090_r = node1084_r & pixel[630];
      node1090_l = node1084_r & ~pixel[630];
      node1091_r = node1090_l & pixel[321];
      node1091_l = node1090_l & ~pixel[321];
      node1092 = node1091_l;
      node1093 = node1091_r;
      node1094 = node1090_r;
      node1095_r = node877_r & pixel[464];
      node1095_l = node877_r & ~pixel[464];
      node1096_r = node1095_l & pixel[516];
      node1096_l = node1095_l & ~pixel[516];
      node1097_r = node1096_l & pixel[431];
      node1097_l = node1096_l & ~pixel[431];
      node1098_r = node1097_l & pixel[436];
      node1098_l = node1097_l & ~pixel[436];
      node1099_r = node1098_l & pixel[372];
      node1099_l = node1098_l & ~pixel[372];
      node1100_r = node1099_l & pixel[300];
      node1100_l = node1099_l & ~pixel[300];
      node1101_r = node1100_l & pixel[205];
      node1101_l = node1100_l & ~pixel[205];
      node1102 = node1101_l;
      node1103 = node1101_r;
      node1104_r = node1100_r & pixel[544];
      node1104_l = node1100_r & ~pixel[544];
      node1105 = node1104_l;
      node1106 = node1104_r;
      node1107_r = node1099_r & pixel[324];
      node1107_l = node1099_r & ~pixel[324];
      node1108_r = node1107_l & pixel[628];
      node1108_l = node1107_l & ~pixel[628];
      node1109 = node1108_l;
      node1110 = node1108_r;
      node1111_r = node1107_r & pixel[583];
      node1111_l = node1107_r & ~pixel[583];
      node1112 = node1111_l;
      node1113 = node1111_r;
      node1114_r = node1098_r & pixel[546];
      node1114_l = node1098_r & ~pixel[546];
      node1115_r = node1114_l & pixel[655];
      node1115_l = node1114_l & ~pixel[655];
      node1116 = node1115_l;
      node1117 = node1115_r;
      node1118 = node1114_r;
      node1119_r = node1097_r & pixel[95];
      node1119_l = node1097_r & ~pixel[95];
      node1120_r = node1119_l & pixel[272];
      node1120_l = node1119_l & ~pixel[272];
      node1121_r = node1120_l & pixel[440];
      node1121_l = node1120_l & ~pixel[440];
      node1122_r = node1121_l & pixel[295];
      node1122_l = node1121_l & ~pixel[295];
      node1123 = node1122_l;
      node1124 = node1122_r;
      node1125_r = node1121_r & pixel[434];
      node1125_l = node1121_r & ~pixel[434];
      node1126 = node1125_l;
      node1127 = node1125_r;
      node1128_r = node1120_r & pixel[346];
      node1128_l = node1120_r & ~pixel[346];
      node1129_r = node1128_l & pixel[622];
      node1129_l = node1128_l & ~pixel[622];
      node1130 = node1129_l;
      node1131 = node1129_r;
      node1132_r = node1128_r & pixel[628];
      node1132_l = node1128_r & ~pixel[628];
      node1133 = node1132_l;
      node1134 = node1132_r;
      node1135 = node1119_r;
      node1136_r = node1096_r & pixel[489];
      node1136_l = node1096_r & ~pixel[489];
      node1137_r = node1136_l & pixel[630];
      node1137_l = node1136_l & ~pixel[630];
      node1138_r = node1137_l & pixel[163];
      node1138_l = node1137_l & ~pixel[163];
      node1139_r = node1138_l & pixel[721];
      node1139_l = node1138_l & ~pixel[721];
      node1140_r = node1139_l & pixel[522];
      node1140_l = node1139_l & ~pixel[522];
      node1141 = node1140_l;
      node1142 = node1140_r;
      node1143 = node1139_r;
      node1144_r = node1138_r & pixel[155];
      node1144_l = node1138_r & ~pixel[155];
      node1145_r = node1144_l & pixel[302];
      node1145_l = node1144_l & ~pixel[302];
      node1146 = node1145_l;
      node1147 = node1145_r;
      node1148 = node1144_r;
      node1149_r = node1137_r & pixel[290];
      node1149_l = node1137_r & ~pixel[290];
      node1150_r = node1149_l & pixel[352];
      node1150_l = node1149_l & ~pixel[352];
      node1151_r = node1150_l & pixel[652];
      node1151_l = node1150_l & ~pixel[652];
      node1152 = node1151_l;
      node1153 = node1151_r;
      node1154_r = node1150_r & pixel[610];
      node1154_l = node1150_r & ~pixel[610];
      node1155 = node1154_l;
      node1156 = node1154_r;
      node1157 = node1149_r;
      node1158_r = node1136_r & pixel[470];
      node1158_l = node1136_r & ~pixel[470];
      node1159_r = node1158_l & pixel[190];
      node1159_l = node1158_l & ~pixel[190];
      node1160_r = node1159_l & pixel[637];
      node1160_l = node1159_l & ~pixel[637];
      node1161_r = node1160_l & pixel[541];
      node1161_l = node1160_l & ~pixel[541];
      node1162 = node1161_l;
      node1163 = node1161_r;
      node1164_r = node1160_r & pixel[182];
      node1164_l = node1160_r & ~pixel[182];
      node1165 = node1164_l;
      node1166 = node1164_r;
      node1167_r = node1159_r & pixel[385];
      node1167_l = node1159_r & ~pixel[385];
      node1168_r = node1167_l & pixel[403];
      node1168_l = node1167_l & ~pixel[403];
      node1169 = node1168_l;
      node1170 = node1168_r;
      node1171 = node1167_r;
      node1172_r = node1158_r & pixel[235];
      node1172_l = node1158_r & ~pixel[235];
      node1173_r = node1172_l & pixel[437];
      node1173_l = node1172_l & ~pixel[437];
      node1174_r = node1173_l & pixel[508];
      node1174_l = node1173_l & ~pixel[508];
      node1175 = node1174_l;
      node1176 = node1174_r;
      node1177 = node1173_r;
      node1178_r = node1172_r & pixel[401];
      node1178_l = node1172_r & ~pixel[401];
      node1179_r = node1178_l & pixel[329];
      node1179_l = node1178_l & ~pixel[329];
      node1180 = node1179_l;
      node1181 = node1179_r;
      node1182_r = node1178_r & pixel[244];
      node1182_l = node1178_r & ~pixel[244];
      node1183 = node1182_l;
      node1184 = node1182_r;
      node1185_r = node1095_r & pixel[349];
      node1185_l = node1095_r & ~pixel[349];
      node1186_r = node1185_l & pixel[316];
      node1186_l = node1185_l & ~pixel[316];
      node1187_r = node1186_l & pixel[293];
      node1187_l = node1186_l & ~pixel[293];
      node1188_r = node1187_l & pixel[690];
      node1188_l = node1187_l & ~pixel[690];
      node1189_r = node1188_l & pixel[631];
      node1189_l = node1188_l & ~pixel[631];
      node1190_r = node1189_l & pixel[284];
      node1190_l = node1189_l & ~pixel[284];
      node1191 = node1190_l;
      node1192 = node1190_r;
      node1193_r = node1189_r & pixel[400];
      node1193_l = node1189_r & ~pixel[400];
      node1194 = node1193_l;
      node1195 = node1193_r;
      node1196_r = node1188_r & pixel[358];
      node1196_l = node1188_r & ~pixel[358];
      node1197_r = node1196_l & pixel[244];
      node1197_l = node1196_l & ~pixel[244];
      node1198 = node1197_l;
      node1199 = node1197_r;
      node1200_r = node1196_r & pixel[570];
      node1200_l = node1196_r & ~pixel[570];
      node1201 = node1200_l;
      node1202 = node1200_r;
      node1203_r = node1187_r & pixel[373];
      node1203_l = node1187_r & ~pixel[373];
      node1204_r = node1203_l & pixel[685];
      node1204_l = node1203_l & ~pixel[685];
      node1205_r = node1204_l & pixel[623];
      node1205_l = node1204_l & ~pixel[623];
      node1206 = node1205_l;
      node1207 = node1205_r;
      node1208 = node1204_r;
      node1209_r = node1203_r & pixel[102];
      node1209_l = node1203_r & ~pixel[102];
      node1210_r = node1209_l & pixel[355];
      node1210_l = node1209_l & ~pixel[355];
      node1211 = node1210_l;
      node1212 = node1210_r;
      node1213_r = node1209_r & pixel[620];
      node1213_l = node1209_r & ~pixel[620];
      node1214 = node1213_l;
      node1215 = node1213_r;
      node1216_r = node1186_r & pixel[570];
      node1216_l = node1186_r & ~pixel[570];
      node1217_r = node1216_l & pixel[580];
      node1217_l = node1216_l & ~pixel[580];
      node1218_r = node1217_l & pixel[625];
      node1218_l = node1217_l & ~pixel[625];
      node1219_r = node1218_l & pixel[579];
      node1219_l = node1218_l & ~pixel[579];
      node1220 = node1219_l;
      node1221 = node1219_r;
      node1222_r = node1218_r & pixel[468];
      node1222_l = node1218_r & ~pixel[468];
      node1223 = node1222_l;
      node1224 = node1222_r;
      node1225_r = node1217_r & pixel[208];
      node1225_l = node1217_r & ~pixel[208];
      node1226_r = node1225_l & pixel[595];
      node1226_l = node1225_l & ~pixel[595];
      node1227 = node1226_l;
      node1228 = node1226_r;
      node1229_r = node1225_r & pixel[355];
      node1229_l = node1225_r & ~pixel[355];
      node1230 = node1229_l;
      node1231 = node1229_r;
      node1232_r = node1216_r & pixel[435];
      node1232_l = node1216_r & ~pixel[435];
      node1233_r = node1232_l & pixel[318];
      node1233_l = node1232_l & ~pixel[318];
      node1234_r = node1233_l & pixel[128];
      node1234_l = node1233_l & ~pixel[128];
      node1235 = node1234_l;
      node1236 = node1234_r;
      node1237_r = node1233_r & pixel[625];
      node1237_l = node1233_r & ~pixel[625];
      node1238 = node1237_l;
      node1239 = node1237_r;
      node1240_r = node1232_r & pixel[214];
      node1240_l = node1232_r & ~pixel[214];
      node1241_r = node1240_l & pixel[357];
      node1241_l = node1240_l & ~pixel[357];
      node1242 = node1241_l;
      node1243 = node1241_r;
      node1244_r = node1240_r & pixel[468];
      node1244_l = node1240_r & ~pixel[468];
      node1245 = node1244_l;
      node1246 = node1244_r;
      node1247_r = node1185_r & pixel[216];
      node1247_l = node1185_r & ~pixel[216];
      node1248_r = node1247_l & pixel[104];
      node1248_l = node1247_l & ~pixel[104];
      node1249_r = node1248_l & pixel[351];
      node1249_l = node1248_l & ~pixel[351];
      node1250_r = node1249_l & pixel[514];
      node1250_l = node1249_l & ~pixel[514];
      node1251_r = node1250_l & pixel[624];
      node1251_l = node1250_l & ~pixel[624];
      node1252 = node1251_l;
      node1253 = node1251_r;
      node1254_r = node1250_r & pixel[654];
      node1254_l = node1250_r & ~pixel[654];
      node1255 = node1254_l;
      node1256 = node1254_r;
      node1257_r = node1249_r & pixel[520];
      node1257_l = node1249_r & ~pixel[520];
      node1258_r = node1257_l & pixel[325];
      node1258_l = node1257_l & ~pixel[325];
      node1259 = node1258_l;
      node1260 = node1258_r;
      node1261_r = node1257_r & pixel[268];
      node1261_l = node1257_r & ~pixel[268];
      node1262 = node1261_l;
      node1263 = node1261_r;
      node1264_r = node1248_r & pixel[242];
      node1264_l = node1248_r & ~pixel[242];
      node1265 = node1264_l;
      node1266_r = node1264_r & pixel[353];
      node1266_l = node1264_r & ~pixel[353];
      node1267 = node1266_l;
      node1268 = node1266_r;
      node1269_r = node1247_r & pixel[272];
      node1269_l = node1247_r & ~pixel[272];
      node1270_r = node1269_l & pixel[331];
      node1270_l = node1269_l & ~pixel[331];
      node1271_r = node1270_l & pixel[514];
      node1271_l = node1270_l & ~pixel[514];
      node1272_r = node1271_l & pixel[542];
      node1272_l = node1271_l & ~pixel[542];
      node1273 = node1272_l;
      node1274 = node1272_r;
      node1275_r = node1271_r & pixel[221];
      node1275_l = node1271_r & ~pixel[221];
      node1276 = node1275_l;
      node1277 = node1275_r;
      node1278_r = node1270_r & pixel[267];
      node1278_l = node1270_r & ~pixel[267];
      node1279 = node1278_l;
      node1280_r = node1278_r & pixel[158];
      node1280_l = node1278_r & ~pixel[158];
      node1281 = node1280_l;
      node1282 = node1280_r;
      node1283_r = node1269_r & pixel[438];
      node1283_l = node1269_r & ~pixel[438];
      node1284_r = node1283_l & pixel[469];
      node1284_l = node1283_l & ~pixel[469];
      node1285_r = node1284_l & pixel[489];
      node1285_l = node1284_l & ~pixel[489];
      node1286 = node1285_l;
      node1287 = node1285_r;
      node1288 = node1284_r;
      node1289_r = node1283_r & pixel[598];
      node1289_l = node1283_r & ~pixel[598];
      node1290_r = node1289_l & pixel[656];
      node1290_l = node1289_l & ~pixel[656];
      node1291 = node1290_l;
      node1292 = node1290_r;
      node1293_r = node1289_r & pixel[461];
      node1293_l = node1289_r & ~pixel[461];
      node1294 = node1293_l;
      node1295 = node1293_r;
      node1296_r = node876_r & pixel[210];
      node1296_l = node876_r & ~pixel[210];
      node1297_r = node1296_l & pixel[153];
      node1297_l = node1296_l & ~pixel[153];
      node1298_r = node1297_l & pixel[95];
      node1298_l = node1297_l & ~pixel[95];
      node1299_r = node1298_l & pixel[119];
      node1299_l = node1298_l & ~pixel[119];
      node1300_r = node1299_l & pixel[624];
      node1300_l = node1299_l & ~pixel[624];
      node1301_r = node1300_l & pixel[400];
      node1301_l = node1300_l & ~pixel[400];
      node1302_r = node1301_l & pixel[377];
      node1302_l = node1301_l & ~pixel[377];
      node1303_r = node1302_l & pixel[160];
      node1303_l = node1302_l & ~pixel[160];
      node1304 = node1303_l;
      node1305 = node1303_r;
      node1306_r = node1302_r & pixel[459];
      node1306_l = node1302_r & ~pixel[459];
      node1307 = node1306_l;
      node1308 = node1306_r;
      node1309_r = node1301_r & pixel[239];
      node1309_l = node1301_r & ~pixel[239];
      node1310_r = node1309_l & pixel[542];
      node1310_l = node1309_l & ~pixel[542];
      node1311 = node1310_l;
      node1312 = node1310_r;
      node1313_r = node1309_r & pixel[156];
      node1313_l = node1309_r & ~pixel[156];
      node1314 = node1313_l;
      node1315 = node1313_r;
      node1316_r = node1300_r & pixel[566];
      node1316_l = node1300_r & ~pixel[566];
      node1317_r = node1316_l & pixel[576];
      node1317_l = node1316_l & ~pixel[576];
      node1318_r = node1317_l & pixel[399];
      node1318_l = node1317_l & ~pixel[399];
      node1319 = node1318_l;
      node1320 = node1318_r;
      node1321_r = node1317_r & pixel[132];
      node1321_l = node1317_r & ~pixel[132];
      node1322 = node1321_l;
      node1323 = node1321_r;
      node1324_r = node1316_r & pixel[513];
      node1324_l = node1316_r & ~pixel[513];
      node1325_r = node1324_l & pixel[356];
      node1325_l = node1324_l & ~pixel[356];
      node1326 = node1325_l;
      node1327 = node1325_r;
      node1328_r = node1324_r & pixel[495];
      node1328_l = node1324_r & ~pixel[495];
      node1329 = node1328_l;
      node1330 = node1328_r;
      node1331_r = node1299_r & pixel[663];
      node1331_l = node1299_r & ~pixel[663];
      node1332_r = node1331_l & pixel[542];
      node1332_l = node1331_l & ~pixel[542];
      node1333_r = node1332_l & pixel[577];
      node1333_l = node1332_l & ~pixel[577];
      node1334 = node1333_l;
      node1335 = node1333_r;
      node1336_r = node1332_r & pixel[209];
      node1336_l = node1332_r & ~pixel[209];
      node1337_r = node1336_l & pixel[238];
      node1337_l = node1336_l & ~pixel[238];
      node1338 = node1337_l;
      node1339 = node1337_r;
      node1340 = node1336_r;
      node1341_r = node1331_r & pixel[655];
      node1341_l = node1331_r & ~pixel[655];
      node1342 = node1341_l;
      node1343_r = node1341_r & pixel[134];
      node1343_l = node1341_r & ~pixel[134];
      node1344 = node1343_l;
      node1345 = node1343_r;
      node1346_r = node1298_r & pixel[155];
      node1346_l = node1298_r & ~pixel[155];
      node1347_r = node1346_l & pixel[130];
      node1347_l = node1346_l & ~pixel[130];
      node1348_r = node1347_l & pixel[547];
      node1348_l = node1347_l & ~pixel[547];
      node1349_r = node1348_l & pixel[267];
      node1349_l = node1348_l & ~pixel[267];
      node1350 = node1349_l;
      node1351 = node1349_r;
      node1352_r = node1348_r & pixel[178];
      node1352_l = node1348_r & ~pixel[178];
      node1353_r = node1352_l & pixel[100];
      node1353_l = node1352_l & ~pixel[100];
      node1354 = node1353_l;
      node1355 = node1353_r;
      node1356 = node1352_r;
      node1357_r = node1347_r & pixel[345];
      node1357_l = node1347_r & ~pixel[345];
      node1358_r = node1357_l & pixel[549];
      node1358_l = node1357_l & ~pixel[549];
      node1359 = node1358_l;
      node1360 = node1358_r;
      node1361 = node1357_r;
      node1362_r = node1346_r & pixel[358];
      node1362_l = node1346_r & ~pixel[358];
      node1363 = node1362_l;
      node1364 = node1362_r;
      node1365_r = node1297_r & pixel[214];
      node1365_l = node1297_r & ~pixel[214];
      node1366_r = node1365_l & pixel[157];
      node1366_l = node1365_l & ~pixel[157];
      node1367_r = node1366_l & pixel[97];
      node1367_l = node1366_l & ~pixel[97];
      node1368_r = node1367_l & pixel[514];
      node1368_l = node1367_l & ~pixel[514];
      node1369_r = node1368_l & pixel[100];
      node1369_l = node1368_l & ~pixel[100];
      node1370_r = node1369_l & pixel[551];
      node1370_l = node1369_l & ~pixel[551];
      node1371 = node1370_l;
      node1372 = node1370_r;
      node1373 = node1369_r;
      node1374_r = node1368_r & pixel[211];
      node1374_l = node1368_r & ~pixel[211];
      node1375_r = node1374_l & pixel[385];
      node1375_l = node1374_l & ~pixel[385];
      node1376 = node1375_l;
      node1377 = node1375_r;
      node1378_r = node1374_r & pixel[538];
      node1378_l = node1374_r & ~pixel[538];
      node1379 = node1378_l;
      node1380 = node1378_r;
      node1381_r = node1367_r & pixel[267];
      node1381_l = node1367_r & ~pixel[267];
      node1382_r = node1381_l & pixel[266];
      node1382_l = node1381_l & ~pixel[266];
      node1383_r = node1382_l & pixel[294];
      node1383_l = node1382_l & ~pixel[294];
      node1384 = node1383_l;
      node1385 = node1383_r;
      node1386 = node1382_r;
      node1387_r = node1381_r & pixel[212];
      node1387_l = node1381_r & ~pixel[212];
      node1388 = node1387_l;
      node1389 = node1387_r;
      node1390_r = node1366_r & pixel[659];
      node1390_l = node1366_r & ~pixel[659];
      node1391_r = node1390_l & pixel[234];
      node1391_l = node1390_l & ~pixel[234];
      node1392_r = node1391_l & pixel[463];
      node1392_l = node1391_l & ~pixel[463];
      node1393_r = node1392_l & pixel[441];
      node1393_l = node1392_l & ~pixel[441];
      node1394 = node1393_l;
      node1395 = node1393_r;
      node1396_r = node1392_r & pixel[612];
      node1396_l = node1392_r & ~pixel[612];
      node1397 = node1396_l;
      node1398 = node1396_r;
      node1399_r = node1391_r & pixel[621];
      node1399_l = node1391_r & ~pixel[621];
      node1400_r = node1399_l & pixel[514];
      node1400_l = node1399_l & ~pixel[514];
      node1401 = node1400_l;
      node1402 = node1400_r;
      node1403_r = node1399_r & pixel[627];
      node1403_l = node1399_r & ~pixel[627];
      node1404 = node1403_l;
      node1405 = node1403_r;
      node1406_r = node1390_r & pixel[131];
      node1406_l = node1390_r & ~pixel[131];
      node1407_r = node1406_l & pixel[345];
      node1407_l = node1406_l & ~pixel[345];
      node1408_r = node1407_l & pixel[510];
      node1408_l = node1407_l & ~pixel[510];
      node1409 = node1408_l;
      node1410 = node1408_r;
      node1411_r = node1407_r & pixel[510];
      node1411_l = node1407_r & ~pixel[510];
      node1412 = node1411_l;
      node1413 = node1411_r;
      node1414_r = node1406_r & pixel[435];
      node1414_l = node1406_r & ~pixel[435];
      node1415_r = node1414_l & pixel[324];
      node1415_l = node1414_l & ~pixel[324];
      node1416 = node1415_l;
      node1417 = node1415_r;
      node1418 = node1414_r;
      node1419_r = node1365_r & pixel[517];
      node1419_l = node1365_r & ~pixel[517];
      node1420_r = node1419_l & pixel[349];
      node1420_l = node1419_l & ~pixel[349];
      node1421_r = node1420_l & pixel[127];
      node1421_l = node1420_l & ~pixel[127];
      node1422_r = node1421_l & pixel[683];
      node1422_l = node1421_l & ~pixel[683];
      node1423_r = node1422_l & pixel[567];
      node1423_l = node1422_l & ~pixel[567];
      node1424 = node1423_l;
      node1425 = node1423_r;
      node1426_r = node1422_r & pixel[327];
      node1426_l = node1422_r & ~pixel[327];
      node1427 = node1426_l;
      node1428 = node1426_r;
      node1429_r = node1421_r & pixel[373];
      node1429_l = node1421_r & ~pixel[373];
      node1430_r = node1429_l & pixel[607];
      node1430_l = node1429_l & ~pixel[607];
      node1431 = node1430_l;
      node1432 = node1430_r;
      node1433_r = node1429_r & pixel[636];
      node1433_l = node1429_r & ~pixel[636];
      node1434 = node1433_l;
      node1435 = node1433_r;
      node1436_r = node1420_r & pixel[264];
      node1436_l = node1420_r & ~pixel[264];
      node1437_r = node1436_l & pixel[317];
      node1437_l = node1436_l & ~pixel[317];
      node1438_r = node1437_l & pixel[468];
      node1438_l = node1437_l & ~pixel[468];
      node1439 = node1438_l;
      node1440 = node1438_r;
      node1441_r = node1437_r & pixel[381];
      node1441_l = node1437_r & ~pixel[381];
      node1442 = node1441_l;
      node1443 = node1441_r;
      node1444_r = node1436_r & pixel[595];
      node1444_l = node1436_r & ~pixel[595];
      node1445_r = node1444_l & pixel[184];
      node1445_l = node1444_l & ~pixel[184];
      node1446 = node1445_l;
      node1447 = node1445_r;
      node1448_r = node1444_r & pixel[665];
      node1448_l = node1444_r & ~pixel[665];
      node1449 = node1448_l;
      node1450 = node1448_r;
      node1451_r = node1419_r & pixel[569];
      node1451_l = node1419_r & ~pixel[569];
      node1452_r = node1451_l & pixel[657];
      node1452_l = node1451_l & ~pixel[657];
      node1453_r = node1452_l & pixel[314];
      node1453_l = node1452_l & ~pixel[314];
      node1454_r = node1453_l & pixel[317];
      node1454_l = node1453_l & ~pixel[317];
      node1455 = node1454_l;
      node1456 = node1454_r;
      node1457 = node1453_r;
      node1458_r = node1452_r & pixel[235];
      node1458_l = node1452_r & ~pixel[235];
      node1459_r = node1458_l & pixel[343];
      node1459_l = node1458_l & ~pixel[343];
      node1460 = node1459_l;
      node1461 = node1459_r;
      node1462_r = node1458_r & pixel[183];
      node1462_l = node1458_r & ~pixel[183];
      node1463 = node1462_l;
      node1464 = node1462_r;
      node1465_r = node1451_r & pixel[430];
      node1465_l = node1451_r & ~pixel[430];
      node1466_r = node1465_l & pixel[404];
      node1466_l = node1465_l & ~pixel[404];
      node1467_r = node1466_l & pixel[344];
      node1467_l = node1466_l & ~pixel[344];
      node1468 = node1467_l;
      node1469 = node1467_r;
      node1470_r = node1466_r & pixel[213];
      node1470_l = node1466_r & ~pixel[213];
      node1471 = node1470_l;
      node1472 = node1470_r;
      node1473_r = node1465_r & pixel[235];
      node1473_l = node1465_r & ~pixel[235];
      node1474 = node1473_l;
      node1475_r = node1473_r & pixel[543];
      node1475_l = node1473_r & ~pixel[543];
      node1476 = node1475_l;
      node1477 = node1475_r;
      node1478_r = node1296_r & pixel[544];
      node1478_l = node1296_r & ~pixel[544];
      node1479_r = node1478_l & pixel[375];
      node1479_l = node1478_l & ~pixel[375];
      node1480_r = node1479_l & pixel[509];
      node1480_l = node1479_l & ~pixel[509];
      node1481_r = node1480_l & pixel[597];
      node1481_l = node1480_l & ~pixel[597];
      node1482_r = node1481_l & pixel[496];
      node1482_l = node1481_l & ~pixel[496];
      node1483_r = node1482_l & pixel[625];
      node1483_l = node1482_l & ~pixel[625];
      node1484_r = node1483_l & pixel[236];
      node1484_l = node1483_l & ~pixel[236];
      node1485 = node1484_l;
      node1486 = node1484_r;
      node1487_r = node1483_r & pixel[545];
      node1487_l = node1483_r & ~pixel[545];
      node1488 = node1487_l;
      node1489 = node1487_r;
      node1490_r = node1482_r & pixel[398];
      node1490_l = node1482_r & ~pixel[398];
      node1491_r = node1490_l & pixel[344];
      node1491_l = node1490_l & ~pixel[344];
      node1492 = node1491_l;
      node1493 = node1491_r;
      node1494_r = node1490_r & pixel[208];
      node1494_l = node1490_r & ~pixel[208];
      node1495 = node1494_l;
      node1496 = node1494_r;
      node1497_r = node1481_r & pixel[433];
      node1497_l = node1481_r & ~pixel[433];
      node1498_r = node1497_l & pixel[321];
      node1498_l = node1497_l & ~pixel[321];
      node1499_r = node1498_l & pixel[212];
      node1499_l = node1498_l & ~pixel[212];
      node1500 = node1499_l;
      node1501 = node1499_r;
      node1502_r = node1498_r & pixel[127];
      node1502_l = node1498_r & ~pixel[127];
      node1503 = node1502_l;
      node1504 = node1502_r;
      node1505_r = node1497_r & pixel[123];
      node1505_l = node1497_r & ~pixel[123];
      node1506_r = node1505_l & pixel[401];
      node1506_l = node1505_l & ~pixel[401];
      node1507 = node1506_l;
      node1508 = node1506_r;
      node1509 = node1505_r;
      node1510_r = node1480_r & pixel[370];
      node1510_l = node1480_r & ~pixel[370];
      node1511_r = node1510_l & pixel[514];
      node1511_l = node1510_l & ~pixel[514];
      node1512_r = node1511_l & pixel[327];
      node1512_l = node1511_l & ~pixel[327];
      node1513_r = node1512_l & pixel[151];
      node1513_l = node1512_l & ~pixel[151];
      node1514 = node1513_l;
      node1515 = node1513_r;
      node1516_r = node1512_r & pixel[434];
      node1516_l = node1512_r & ~pixel[434];
      node1517 = node1516_l;
      node1518 = node1516_r;
      node1519_r = node1511_r & pixel[320];
      node1519_l = node1511_r & ~pixel[320];
      node1520_r = node1519_l & pixel[628];
      node1520_l = node1519_l & ~pixel[628];
      node1521 = node1520_l;
      node1522 = node1520_r;
      node1523_r = node1519_r & pixel[274];
      node1523_l = node1519_r & ~pixel[274];
      node1524 = node1523_l;
      node1525 = node1523_r;
      node1526_r = node1510_r & pixel[598];
      node1526_l = node1510_r & ~pixel[598];
      node1527_r = node1526_l & pixel[266];
      node1527_l = node1526_l & ~pixel[266];
      node1528_r = node1527_l & pixel[599];
      node1528_l = node1527_l & ~pixel[599];
      node1529 = node1528_l;
      node1530 = node1528_r;
      node1531_r = node1527_r & pixel[122];
      node1531_l = node1527_r & ~pixel[122];
      node1532 = node1531_l;
      node1533 = node1531_r;
      node1534 = node1526_r;
      node1535_r = node1479_r & pixel[274];
      node1535_l = node1479_r & ~pixel[274];
      node1536_r = node1535_l & pixel[513];
      node1536_l = node1535_l & ~pixel[513];
      node1537_r = node1536_l & pixel[188];
      node1537_l = node1536_l & ~pixel[188];
      node1538_r = node1537_l & pixel[598];
      node1538_l = node1537_l & ~pixel[598];
      node1539_r = node1538_l & pixel[203];
      node1539_l = node1538_l & ~pixel[203];
      node1540 = node1539_l;
      node1541 = node1539_r;
      node1542_r = node1538_r & pixel[431];
      node1542_l = node1538_r & ~pixel[431];
      node1543 = node1542_l;
      node1544 = node1542_r;
      node1545_r = node1537_r & pixel[372];
      node1545_l = node1537_r & ~pixel[372];
      node1546_r = node1545_l & pixel[184];
      node1546_l = node1545_l & ~pixel[184];
      node1547 = node1546_l;
      node1548 = node1546_r;
      node1549_r = node1545_r & pixel[213];
      node1549_l = node1545_r & ~pixel[213];
      node1550 = node1549_l;
      node1551 = node1549_r;
      node1552_r = node1536_r & pixel[299];
      node1552_l = node1536_r & ~pixel[299];
      node1553_r = node1552_l & pixel[270];
      node1553_l = node1552_l & ~pixel[270];
      node1554_r = node1553_l & pixel[574];
      node1554_l = node1553_l & ~pixel[574];
      node1555 = node1554_l;
      node1556 = node1554_r;
      node1557_r = node1553_r & pixel[490];
      node1557_l = node1553_r & ~pixel[490];
      node1558 = node1557_l;
      node1559 = node1557_r;
      node1560_r = node1552_r & pixel[712];
      node1560_l = node1552_r & ~pixel[712];
      node1561_r = node1560_l & pixel[626];
      node1561_l = node1560_l & ~pixel[626];
      node1562 = node1561_l;
      node1563 = node1561_r;
      node1564_r = node1560_r & pixel[568];
      node1564_l = node1560_r & ~pixel[568];
      node1565 = node1564_l;
      node1566 = node1564_r;
      node1567_r = node1535_r & pixel[397];
      node1567_l = node1535_r & ~pixel[397];
      node1568_r = node1567_l & pixel[512];
      node1568_l = node1567_l & ~pixel[512];
      node1569_r = node1568_l & pixel[481];
      node1569_l = node1568_l & ~pixel[481];
      node1570_r = node1569_l & pixel[212];
      node1570_l = node1569_l & ~pixel[212];
      node1571 = node1570_l;
      node1572 = node1570_r;
      node1573_r = node1569_r & pixel[149];
      node1573_l = node1569_r & ~pixel[149];
      node1574 = node1573_l;
      node1575 = node1573_r;
      node1576_r = node1568_r & pixel[372];
      node1576_l = node1568_r & ~pixel[372];
      node1577_r = node1576_l & pixel[236];
      node1577_l = node1576_l & ~pixel[236];
      node1578 = node1577_l;
      node1579 = node1577_r;
      node1580_r = node1576_r & pixel[432];
      node1580_l = node1576_r & ~pixel[432];
      node1581 = node1580_l;
      node1582 = node1580_r;
      node1583_r = node1567_r & pixel[387];
      node1583_l = node1567_r & ~pixel[387];
      node1584_r = node1583_l & pixel[576];
      node1584_l = node1583_l & ~pixel[576];
      node1585_r = node1584_l & pixel[488];
      node1585_l = node1584_l & ~pixel[488];
      node1586 = node1585_l;
      node1587 = node1585_r;
      node1588_r = node1584_r & pixel[577];
      node1588_l = node1584_r & ~pixel[577];
      node1589 = node1588_l;
      node1590 = node1588_r;
      node1591_r = node1583_r & pixel[487];
      node1591_l = node1583_r & ~pixel[487];
      node1592 = node1591_l;
      node1593 = node1591_r;
      node1594_r = node1478_r & pixel[290];
      node1594_l = node1478_r & ~pixel[290];
      node1595_r = node1594_l & pixel[320];
      node1595_l = node1594_l & ~pixel[320];
      node1596_r = node1595_l & pixel[655];
      node1596_l = node1595_l & ~pixel[655];
      node1597_r = node1596_l & pixel[661];
      node1597_l = node1596_l & ~pixel[661];
      node1598_r = node1597_l & pixel[248];
      node1598_l = node1597_l & ~pixel[248];
      node1599_r = node1598_l & pixel[316];
      node1599_l = node1598_l & ~pixel[316];
      node1600 = node1599_l;
      node1601 = node1599_r;
      node1602_r = node1598_r & pixel[324];
      node1602_l = node1598_r & ~pixel[324];
      node1603 = node1602_l;
      node1604 = node1602_r;
      node1605_r = node1597_r & pixel[128];
      node1605_l = node1597_r & ~pixel[128];
      node1606_r = node1605_l & pixel[343];
      node1606_l = node1605_l & ~pixel[343];
      node1607 = node1606_l;
      node1608 = node1606_r;
      node1609 = node1605_r;
      node1610_r = node1596_r & pixel[710];
      node1610_l = node1596_r & ~pixel[710];
      node1611_r = node1610_l & pixel[487];
      node1611_l = node1610_l & ~pixel[487];
      node1612_r = node1611_l & pixel[302];
      node1612_l = node1611_l & ~pixel[302];
      node1613 = node1612_l;
      node1614 = node1612_r;
      node1615_r = node1611_r & pixel[549];
      node1615_l = node1611_r & ~pixel[549];
      node1616 = node1615_l;
      node1617 = node1615_r;
      node1618_r = node1610_r & pixel[435];
      node1618_l = node1610_r & ~pixel[435];
      node1619 = node1618_l;
      node1620 = node1618_r;
      node1621_r = node1595_r & pixel[655];
      node1621_l = node1595_r & ~pixel[655];
      node1622_r = node1621_l & pixel[234];
      node1622_l = node1621_l & ~pixel[234];
      node1623_r = node1622_l & pixel[271];
      node1623_l = node1622_l & ~pixel[271];
      node1624_r = node1623_l & pixel[541];
      node1624_l = node1623_l & ~pixel[541];
      node1625 = node1624_l;
      node1626 = node1624_r;
      node1627_r = node1623_r & pixel[319];
      node1627_l = node1623_r & ~pixel[319];
      node1628 = node1627_l;
      node1629 = node1627_r;
      node1630_r = node1622_r & pixel[431];
      node1630_l = node1622_r & ~pixel[431];
      node1631 = node1630_l;
      node1632_r = node1630_r & pixel[518];
      node1632_l = node1630_r & ~pixel[518];
      node1633 = node1632_l;
      node1634 = node1632_r;
      node1635_r = node1621_r & pixel[659];
      node1635_l = node1621_r & ~pixel[659];
      node1636_r = node1635_l & pixel[241];
      node1636_l = node1635_l & ~pixel[241];
      node1637_r = node1636_l & pixel[596];
      node1637_l = node1636_l & ~pixel[596];
      node1638 = node1637_l;
      node1639 = node1637_r;
      node1640_r = node1636_r & pixel[625];
      node1640_l = node1636_r & ~pixel[625];
      node1641 = node1640_l;
      node1642 = node1640_r;
      node1643_r = node1635_r & pixel[665];
      node1643_l = node1635_r & ~pixel[665];
      node1644_r = node1643_l & pixel[439];
      node1644_l = node1643_l & ~pixel[439];
      node1645 = node1644_l;
      node1646 = node1644_r;
      node1647 = node1643_r;
      node1648_r = node1594_r & pixel[578];
      node1648_l = node1594_r & ~pixel[578];
      node1649_r = node1648_l & pixel[127];
      node1649_l = node1648_l & ~pixel[127];
      node1650_r = node1649_l & pixel[213];
      node1650_l = node1649_l & ~pixel[213];
      node1651_r = node1650_l & pixel[177];
      node1651_l = node1650_l & ~pixel[177];
      node1652_r = node1651_l & pixel[552];
      node1652_l = node1651_l & ~pixel[552];
      node1653 = node1652_l;
      node1654 = node1652_r;
      node1655_r = node1651_r & pixel[466];
      node1655_l = node1651_r & ~pixel[466];
      node1656 = node1655_l;
      node1657 = node1655_r;
      node1658_r = node1650_r & pixel[511];
      node1658_l = node1650_r & ~pixel[511];
      node1659_r = node1658_l & pixel[300];
      node1659_l = node1658_l & ~pixel[300];
      node1660 = node1659_l;
      node1661 = node1659_r;
      node1662_r = node1658_r & pixel[105];
      node1662_l = node1658_r & ~pixel[105];
      node1663 = node1662_l;
      node1664 = node1662_r;
      node1665_r = node1649_r & pixel[318];
      node1665_l = node1649_r & ~pixel[318];
      node1666_r = node1665_l & pixel[330];
      node1666_l = node1665_l & ~pixel[330];
      node1667_r = node1666_l & pixel[549];
      node1667_l = node1666_l & ~pixel[549];
      node1668 = node1667_l;
      node1669 = node1667_r;
      node1670 = node1666_r;
      node1671_r = node1665_r & pixel[205];
      node1671_l = node1665_r & ~pixel[205];
      node1672_r = node1671_l & pixel[188];
      node1672_l = node1671_l & ~pixel[188];
      node1673 = node1672_l;
      node1674 = node1672_r;
      node1675 = node1671_r;
      node1676_r = node1648_r & pixel[99];
      node1676_l = node1648_r & ~pixel[99];
      node1677_r = node1676_l & pixel[130];
      node1677_l = node1676_l & ~pixel[130];
      node1678_r = node1677_l & pixel[658];
      node1678_l = node1677_l & ~pixel[658];
      node1679_r = node1678_l & pixel[528];
      node1679_l = node1678_l & ~pixel[528];
      node1680 = node1679_l;
      node1681 = node1679_r;
      node1682_r = node1678_r & pixel[461];
      node1682_l = node1678_r & ~pixel[461];
      node1683 = node1682_l;
      node1684 = node1682_r;
      node1685_r = node1677_r & pixel[188];
      node1685_l = node1677_r & ~pixel[188];
      node1686_r = node1685_l & pixel[178];
      node1686_l = node1685_l & ~pixel[178];
      node1687 = node1686_l;
      node1688 = node1686_r;
      node1689_r = node1685_r & pixel[300];
      node1689_l = node1685_r & ~pixel[300];
      node1690 = node1689_l;
      node1691 = node1689_r;
      node1692_r = node1676_r & pixel[214];
      node1692_l = node1676_r & ~pixel[214];
      node1693_r = node1692_l & pixel[94];
      node1693_l = node1692_l & ~pixel[94];
      node1694_r = node1693_l & pixel[512];
      node1694_l = node1693_l & ~pixel[512];
      node1695 = node1694_l;
      node1696 = node1694_r;
      node1697_r = node1693_r & pixel[185];
      node1697_l = node1693_r & ~pixel[185];
      node1698 = node1697_l;
      node1699 = node1697_r;
      node1700_r = node1692_r & pixel[439];
      node1700_l = node1692_r & ~pixel[439];
      node1701_r = node1700_l & pixel[270];
      node1701_l = node1700_l & ~pixel[270];
      node1702 = node1701_l;
      node1703 = node1701_r;
      node1704_r = node1700_r & pixel[490];
      node1704_l = node1700_r & ~pixel[490];
      node1705 = node1704_l;
      node1706 = node1704_r;
      result0 = node80 | node95 | node105 | node119 | node122 | node135 | node144 | node145 | node157 | node174 | node281 | node417 | node432 | node457 | node465 | node473 | node493 | node523 | node524 | node529 | node530 | node560 | node575 | node578 | node620 | node806 | node885 | node903 | node904 | node908 | node917 | node932 | node937 | node939 | node947 | node950 | node953 | node968 | node980 | node993 | node1024 | node1033 | node1040 | node1046 | node1049 | node1050 | node1061 | node1062 | node1073 | node1078 | node1082 | node1087 | node1102 | node1105 | node1106 | node1109 | node1110 | node1112 | node1113 | node1118 | node1123 | node1126 | node1131 | node1133 | node1134 | node1142 | node1152 | node1153 | node1157 | node1175 | node1181 | node1183 | node1184 | node1212 | node1215 | node1224 | node1238 | node1239 | node1253 | node1256 | node1268 | node1281 | node1282 | node1288 | node1292 | node1294 | node1295 | node1339 | node1386 | node1416 | node1434 | node1469 | node1501 | node1534 | node1566 | node1581 | node1592 | node1614 | node1683 | node1705;
      result1 = node20 | node21 | node181 | node236 | node239 | node240 | node244 | node343 | node582 | node656 | node671 | node1162;
      result2 = node45 | node74 | node76 | node84 | node138 | node167 | node232 | node237 | node245 | node251 | node252 | node254 | node294 | node301 | node305 | node308 | node316 | node320 | node322 | node323 | node326 | node331 | node334 | node335 | node350 | node362 | node370 | node371 | node390 | node399 | node400 | node402 | node406 | node407 | node409 | node416 | node422 | node437 | node444 | node471 | node515 | node556 | node561 | node577 | node585 | node589 | node592 | node641 | node648 | node679 | node691 | node807 | node812 | node818 | node867 | node872 | node889 | node916 | node919 | node926 | node930 | node936 | node940 | node946 | node965 | node969 | node971 | node981 | node1007 | node1009 | node1025 | node1041 | node1047 | node1072 | node1124 | node1130 | node1135 | node1141 | node1156 | node1163 | node1171 | node1176 | node1180 | node1191 | node1194 | node1195 | node1206 | node1207 | node1228 | node1246 | node1263 | node1279 | node1340 | node1355 | node1360 | node1363 | node1380 | node1389 | node1395 | node1397 | node1404 | node1431 | node1432 | node1442 | node1455 | node1468 | node1474 | node1476 | node1477 | node1492 | node1509 | node1521 | node1522 | node1524 | node1575 | node1587 | node1600 | node1607 | node1609 | node1617 | node1628 | node1634 | node1647 | node1657 | node1663 | node1668 | node1669 | node1674 | node1675 | node1681 | node1688 | node1691 | node1703;
      result3 = node10 | node11 | node48 | node66 | node73 | node77 | node89 | node92 | node120 | node126 | node127 | node130 | node137 | node142 | node150 | node151 | node158 | node159 | node163 | node164 | node166 | node170 | node171 | node187 | node188 | node196 | node203 | node210 | node276 | node290 | node312 | node330 | node333 | node351 | node355 | node358 | node368 | node383 | node393 | node448 | node468 | node482 | node486 | node519 | node568 | node571 | node630 | node672 | node675 | node685 | node736 | node775 | node819 | node822 | node826 | node836 | node844 | node864 | node871 | node972 | node1103 | node1148 | node1155 | node1260 | node1394 | node1409 | node1427 | node1439 | node1440 | node1460 | node1488 | node1504 | node1517 | node1541 | node1544 | node1548 | node1572 | node1613 | node1631 | node1633 | node1645 | node1646 | node1699;
      result4 = node36 | node41 | node219 | node265 | node342 | node356 | node377 | node378 | node415 | node522 | node562 | node600 | node627 | node640 | node708 | node711 | node723 | node740 | node757 | node833 | node834 | node837 | node888 | node911 | node962 | node964 | node977 | node988 | node994 | node998 | node1065 | node1116 | node1165 | node1192 | node1198 | node1227 | node1291 | node1304 | node1305 | node1311 | node1312 | node1315 | node1319 | node1320 | node1334 | node1342 | node1361 | node1371 | node1424 | node1446 | node1450 | node1456 | node1457 | node1463 | node1495 | node1529 | node1533 | node1547 | node1550 | node1559 | node1562 | node1571 | node1589 | node1625 | node1629 | node1638 | node1641 | node1653;
      result5 = node13 | node18 | node35 | node44 | node57 | node91 | node98 | node99 | node102 | node106 | node107 | node111 | node129 | node134 | node141 | node173 | node184 | node189 | node212 | node260 | node268 | node274 | node283 | node347 | node359 | node382 | node440 | node458 | node460 | node464 | node467 | node479 | node481 | node485 | node488 | node489 | node494 | node495 | node496 | node503 | node509 | node511 | node516 | node518 | node533 | node546 | node553 | node554 | node567 | node570 | node615 | node619 | node622 | node632 | node644 | node655 | node684 | node701 | node717 | node732 | node733 | node735 | node738 | node745 | node746 | node748 | node758 | node760 | node764 | node765 | node768 | node772 | node776 | node779 | node788 | node803 | node809 | node841 | node856 | node859 | node874 | node892 | node900 | node901 | node1016 | node1021 | node1027 | node1034 | node1036 | node1037 | node1042 | node1127 | node1146 | node1169 | node1170 | node1199 | node1211 | node1223 | node1230 | node1245 | node1273 | node1277 | node1287 | node1307 | node1322 | node1326 | node1344 | node1351 | node1410 | node1412 | node1417 | node1503 | node1514 | node1543 | node1551 | node1555 | node1604;
      result6 = node14 | node17 | node32 | node33 | node42 | node51 | node81 | node83 | node88 | node229 | node262 | node273 | node277 | node280 | node325 | node348 | node374 | node430 | node438 | node441 | node472 | node510 | node593 | node601 | node625 | node631 | node663 | node665 | node680 | node704 | node712 | node886 | node896 | node920 | node923 | node924 | node927 | node933 | node949 | node954 | node956 | node957 | node961 | node978 | node985 | node987 | node992 | node996 | node999 | node1089 | node1177 | node1214 | node1236 | node1242 | node1243 | node1252 | node1255 | node1265 | node1267 | node1274 | node1276 | node1308 | node1323 | node1330 | node1335 | node1338 | node1350 | node1354 | node1356 | node1359 | node1364 | node1373 | node1376 | node1377 | node1384 | node1385 | node1388 | node1398 | node1401 | node1402 | node1472 | node1500 | node1556 | node1601 | node1626 | node1664 | node1673 | node1687 | node1690 | node1695 | node1696 | node1698 | node1702 | node1706;
      result7 = node25 | node26 | node56 | node59 | node112 | node123 | node154 | node183 | node193 | node201 | node204 | node216 | node217 | node291 | node293 | node297 | node306 | node461 | node478 | node502 | node505 | node506 | node531 | node532 | node540 | node541 | node543 | node544 | node548 | node549 | node574 | node583 | node604 | node605 | node608 | node616 | node647 | node650 | node658 | node666 | node850 | node895 | node907 | node984 | node1014 | node1022 | node1052 | node1060 | node1083 | node1093 | node1603 | node1620;
      result8 = node29 | node64 | node96 | node109 | node153 | node208 | node221 | node230 | node233 | node247 | node248 | node255 | node261 | node269 | node284 | node298 | node300 | node309 | node313 | node315 | node344 | node363 | node364 | node375 | node385 | node392 | node403 | node410 | node423 | node425 | node426 | node429 | node433 | node445 | node447 | node612 | node613 | node623 | node659 | node662 | node674 | node678 | node687 | node688 | node692 | node694 | node695 | node709 | node726 | node727 | node741 | node749 | node750 | node761 | node767 | node773 | node780 | node782 | node783 | node791 | node792 | node795 | node799 | node804 | node811 | node821 | node825 | node828 | node829 | node840 | node843 | node857 | node860 | node865 | node868 | node875 | node1068 | node1071 | node1088 | node1094 | node1117 | node1147 | node1202 | node1208 | node1259 | node1262 | node1286 | node1327 | node1329 | node1345 | node1379 | node1405 | node1413 | node1418 | node1428 | node1435 | node1443 | node1447 | node1449 | node1461 | node1471 | node1489 | node1507 | node1508 | node1515 | node1518 | node1525 | node1558 | node1563 | node1574 | node1578 | node1579 | node1582 | node1586 | node1593 | node1616 | node1639 | node1642 | node1654 | node1656 | node1670 | node1684;
      result9 = node28 | node49 | node52 | node60 | node63 | node67 | node180 | node194 | node197 | node200 | node211 | node220 | node266 | node386 | node389 | node412 | node557 | node586 | node590 | node599 | node607 | node643 | node651 | node702 | node705 | node716 | node719 | node720 | node724 | node789 | node796 | node798 | node849 | node852 | node853 | node893 | node910 | node1006 | node1010 | node1013 | node1017 | node1028 | node1053 | node1059 | node1067 | node1079 | node1081 | node1092 | node1143 | node1166 | node1201 | node1220 | node1221 | node1231 | node1235 | node1314 | node1372 | node1425 | node1464 | node1485 | node1486 | node1493 | node1496 | node1530 | node1532 | node1540 | node1565 | node1590 | node1608 | node1619 | node1660 | node1661 | node1680;

      tree_2 = {result9, result8, result7, result6, result5, result4, result3, result2, result1, result0};
    end
  endfunction

  function [9:0] tree_3;
    input [783:0] pixel;

    reg node0_r;
    reg node0_l;
    reg node1_r;
    reg node1_l;
    reg node2_r;
    reg node2_l;
    reg node3_r;
    reg node3_l;
    reg node4_r;
    reg node4_l;
    reg node5_r;
    reg node5_l;
    reg node6_r;
    reg node6_l;
    reg node7_r;
    reg node7_l;
    reg node8_r;
    reg node8_l;
    reg node9_r;
    reg node9_l;
    reg node10;
    reg node11;
    reg node12_r;
    reg node12_l;
    reg node13;
    reg node14;
    reg node15_r;
    reg node15_l;
    reg node16_r;
    reg node16_l;
    reg node17;
    reg node18;
    reg node19_r;
    reg node19_l;
    reg node20;
    reg node21;
    reg node22_r;
    reg node22_l;
    reg node23_r;
    reg node23_l;
    reg node24_r;
    reg node24_l;
    reg node25;
    reg node26;
    reg node27_r;
    reg node27_l;
    reg node28;
    reg node29;
    reg node30_r;
    reg node30_l;
    reg node31_r;
    reg node31_l;
    reg node32;
    reg node33;
    reg node34_r;
    reg node34_l;
    reg node35;
    reg node36;
    reg node37_r;
    reg node37_l;
    reg node38_r;
    reg node38_l;
    reg node39_r;
    reg node39_l;
    reg node40_r;
    reg node40_l;
    reg node41;
    reg node42;
    reg node43_r;
    reg node43_l;
    reg node44;
    reg node45;
    reg node46_r;
    reg node46_l;
    reg node47_r;
    reg node47_l;
    reg node48;
    reg node49;
    reg node50_r;
    reg node50_l;
    reg node51;
    reg node52;
    reg node53_r;
    reg node53_l;
    reg node54_r;
    reg node54_l;
    reg node55;
    reg node56;
    reg node57_r;
    reg node57_l;
    reg node58;
    reg node59_r;
    reg node59_l;
    reg node60;
    reg node61;
    reg node62_r;
    reg node62_l;
    reg node63_r;
    reg node63_l;
    reg node64_r;
    reg node64_l;
    reg node65_r;
    reg node65_l;
    reg node66_r;
    reg node66_l;
    reg node67;
    reg node68;
    reg node69_r;
    reg node69_l;
    reg node70;
    reg node71;
    reg node72_r;
    reg node72_l;
    reg node73_r;
    reg node73_l;
    reg node74;
    reg node75;
    reg node76_r;
    reg node76_l;
    reg node77;
    reg node78;
    reg node79_r;
    reg node79_l;
    reg node80_r;
    reg node80_l;
    reg node81_r;
    reg node81_l;
    reg node82;
    reg node83;
    reg node84_r;
    reg node84_l;
    reg node85;
    reg node86;
    reg node87_r;
    reg node87_l;
    reg node88_r;
    reg node88_l;
    reg node89;
    reg node90;
    reg node91_r;
    reg node91_l;
    reg node92;
    reg node93;
    reg node94_r;
    reg node94_l;
    reg node95_r;
    reg node95_l;
    reg node96_r;
    reg node96_l;
    reg node97_r;
    reg node97_l;
    reg node98;
    reg node99;
    reg node100_r;
    reg node100_l;
    reg node101;
    reg node102;
    reg node103;
    reg node104_r;
    reg node104_l;
    reg node105_r;
    reg node105_l;
    reg node106_r;
    reg node106_l;
    reg node107;
    reg node108;
    reg node109_r;
    reg node109_l;
    reg node110;
    reg node111;
    reg node112;
    reg node113_r;
    reg node113_l;
    reg node114_r;
    reg node114_l;
    reg node115_r;
    reg node115_l;
    reg node116_r;
    reg node116_l;
    reg node117_r;
    reg node117_l;
    reg node118_r;
    reg node118_l;
    reg node119;
    reg node120;
    reg node121_r;
    reg node121_l;
    reg node122;
    reg node123;
    reg node124_r;
    reg node124_l;
    reg node125_r;
    reg node125_l;
    reg node126;
    reg node127;
    reg node128_r;
    reg node128_l;
    reg node129;
    reg node130;
    reg node131_r;
    reg node131_l;
    reg node132_r;
    reg node132_l;
    reg node133_r;
    reg node133_l;
    reg node134;
    reg node135;
    reg node136_r;
    reg node136_l;
    reg node137;
    reg node138;
    reg node139_r;
    reg node139_l;
    reg node140_r;
    reg node140_l;
    reg node141;
    reg node142;
    reg node143_r;
    reg node143_l;
    reg node144;
    reg node145;
    reg node146_r;
    reg node146_l;
    reg node147_r;
    reg node147_l;
    reg node148_r;
    reg node148_l;
    reg node149_r;
    reg node149_l;
    reg node150;
    reg node151;
    reg node152_r;
    reg node152_l;
    reg node153;
    reg node154;
    reg node155_r;
    reg node155_l;
    reg node156_r;
    reg node156_l;
    reg node157;
    reg node158;
    reg node159_r;
    reg node159_l;
    reg node160;
    reg node161;
    reg node162_r;
    reg node162_l;
    reg node163;
    reg node164_r;
    reg node164_l;
    reg node165;
    reg node166_r;
    reg node166_l;
    reg node167;
    reg node168;
    reg node169_r;
    reg node169_l;
    reg node170_r;
    reg node170_l;
    reg node171_r;
    reg node171_l;
    reg node172_r;
    reg node172_l;
    reg node173_r;
    reg node173_l;
    reg node174;
    reg node175;
    reg node176_r;
    reg node176_l;
    reg node177;
    reg node178;
    reg node179_r;
    reg node179_l;
    reg node180_r;
    reg node180_l;
    reg node181;
    reg node182;
    reg node183_r;
    reg node183_l;
    reg node184;
    reg node185;
    reg node186_r;
    reg node186_l;
    reg node187_r;
    reg node187_l;
    reg node188_r;
    reg node188_l;
    reg node189;
    reg node190;
    reg node191_r;
    reg node191_l;
    reg node192;
    reg node193;
    reg node194_r;
    reg node194_l;
    reg node195_r;
    reg node195_l;
    reg node196;
    reg node197;
    reg node198_r;
    reg node198_l;
    reg node199;
    reg node200;
    reg node201_r;
    reg node201_l;
    reg node202_r;
    reg node202_l;
    reg node203_r;
    reg node203_l;
    reg node204;
    reg node205_r;
    reg node205_l;
    reg node206;
    reg node207;
    reg node208;
    reg node209_r;
    reg node209_l;
    reg node210_r;
    reg node210_l;
    reg node211;
    reg node212;
    reg node213_r;
    reg node213_l;
    reg node214_r;
    reg node214_l;
    reg node215;
    reg node216;
    reg node217;
    reg node218_r;
    reg node218_l;
    reg node219_r;
    reg node219_l;
    reg node220_r;
    reg node220_l;
    reg node221_r;
    reg node221_l;
    reg node222_r;
    reg node222_l;
    reg node223_r;
    reg node223_l;
    reg node224_r;
    reg node224_l;
    reg node225;
    reg node226;
    reg node227_r;
    reg node227_l;
    reg node228;
    reg node229;
    reg node230_r;
    reg node230_l;
    reg node231_r;
    reg node231_l;
    reg node232;
    reg node233;
    reg node234_r;
    reg node234_l;
    reg node235;
    reg node236;
    reg node237_r;
    reg node237_l;
    reg node238_r;
    reg node238_l;
    reg node239_r;
    reg node239_l;
    reg node240;
    reg node241;
    reg node242_r;
    reg node242_l;
    reg node243;
    reg node244;
    reg node245_r;
    reg node245_l;
    reg node246_r;
    reg node246_l;
    reg node247;
    reg node248;
    reg node249_r;
    reg node249_l;
    reg node250;
    reg node251;
    reg node252;
    reg node253_r;
    reg node253_l;
    reg node254_r;
    reg node254_l;
    reg node255_r;
    reg node255_l;
    reg node256_r;
    reg node256_l;
    reg node257_r;
    reg node257_l;
    reg node258;
    reg node259;
    reg node260_r;
    reg node260_l;
    reg node261;
    reg node262;
    reg node263_r;
    reg node263_l;
    reg node264_r;
    reg node264_l;
    reg node265;
    reg node266;
    reg node267_r;
    reg node267_l;
    reg node268;
    reg node269;
    reg node270_r;
    reg node270_l;
    reg node271_r;
    reg node271_l;
    reg node272_r;
    reg node272_l;
    reg node273;
    reg node274;
    reg node275_r;
    reg node275_l;
    reg node276;
    reg node277;
    reg node278_r;
    reg node278_l;
    reg node279_r;
    reg node279_l;
    reg node280;
    reg node281;
    reg node282_r;
    reg node282_l;
    reg node283;
    reg node284;
    reg node285_r;
    reg node285_l;
    reg node286_r;
    reg node286_l;
    reg node287_r;
    reg node287_l;
    reg node288_r;
    reg node288_l;
    reg node289;
    reg node290;
    reg node291_r;
    reg node291_l;
    reg node292;
    reg node293;
    reg node294_r;
    reg node294_l;
    reg node295_r;
    reg node295_l;
    reg node296;
    reg node297;
    reg node298_r;
    reg node298_l;
    reg node299;
    reg node300;
    reg node301_r;
    reg node301_l;
    reg node302_r;
    reg node302_l;
    reg node303_r;
    reg node303_l;
    reg node304;
    reg node305;
    reg node306_r;
    reg node306_l;
    reg node307;
    reg node308;
    reg node309_r;
    reg node309_l;
    reg node310_r;
    reg node310_l;
    reg node311;
    reg node312;
    reg node313;
    reg node314_r;
    reg node314_l;
    reg node315_r;
    reg node315_l;
    reg node316_r;
    reg node316_l;
    reg node317_r;
    reg node317_l;
    reg node318_r;
    reg node318_l;
    reg node319_r;
    reg node319_l;
    reg node320;
    reg node321;
    reg node322_r;
    reg node322_l;
    reg node323;
    reg node324;
    reg node325_r;
    reg node325_l;
    reg node326;
    reg node327_r;
    reg node327_l;
    reg node328;
    reg node329;
    reg node330;
    reg node331_r;
    reg node331_l;
    reg node332_r;
    reg node332_l;
    reg node333_r;
    reg node333_l;
    reg node334_r;
    reg node334_l;
    reg node335;
    reg node336;
    reg node337;
    reg node338;
    reg node339_r;
    reg node339_l;
    reg node340_r;
    reg node340_l;
    reg node341_r;
    reg node341_l;
    reg node342;
    reg node343;
    reg node344;
    reg node345_r;
    reg node345_l;
    reg node346;
    reg node347;
    reg node348_r;
    reg node348_l;
    reg node349_r;
    reg node349_l;
    reg node350_r;
    reg node350_l;
    reg node351;
    reg node352;
    reg node353;
    reg node354_r;
    reg node354_l;
    reg node355;
    reg node356;
    reg node357_r;
    reg node357_l;
    reg node358_r;
    reg node358_l;
    reg node359_r;
    reg node359_l;
    reg node360_r;
    reg node360_l;
    reg node361_r;
    reg node361_l;
    reg node362_r;
    reg node362_l;
    reg node363_r;
    reg node363_l;
    reg node364_r;
    reg node364_l;
    reg node365;
    reg node366;
    reg node367_r;
    reg node367_l;
    reg node368;
    reg node369;
    reg node370_r;
    reg node370_l;
    reg node371_r;
    reg node371_l;
    reg node372;
    reg node373;
    reg node374_r;
    reg node374_l;
    reg node375;
    reg node376;
    reg node377_r;
    reg node377_l;
    reg node378_r;
    reg node378_l;
    reg node379_r;
    reg node379_l;
    reg node380;
    reg node381;
    reg node382_r;
    reg node382_l;
    reg node383;
    reg node384;
    reg node385_r;
    reg node385_l;
    reg node386_r;
    reg node386_l;
    reg node387;
    reg node388;
    reg node389_r;
    reg node389_l;
    reg node390;
    reg node391;
    reg node392_r;
    reg node392_l;
    reg node393_r;
    reg node393_l;
    reg node394_r;
    reg node394_l;
    reg node395_r;
    reg node395_l;
    reg node396;
    reg node397;
    reg node398_r;
    reg node398_l;
    reg node399;
    reg node400;
    reg node401_r;
    reg node401_l;
    reg node402_r;
    reg node402_l;
    reg node403;
    reg node404;
    reg node405_r;
    reg node405_l;
    reg node406;
    reg node407;
    reg node408;
    reg node409_r;
    reg node409_l;
    reg node410_r;
    reg node410_l;
    reg node411_r;
    reg node411_l;
    reg node412_r;
    reg node412_l;
    reg node413_r;
    reg node413_l;
    reg node414;
    reg node415;
    reg node416_r;
    reg node416_l;
    reg node417;
    reg node418;
    reg node419_r;
    reg node419_l;
    reg node420_r;
    reg node420_l;
    reg node421;
    reg node422;
    reg node423_r;
    reg node423_l;
    reg node424;
    reg node425;
    reg node426_r;
    reg node426_l;
    reg node427;
    reg node428_r;
    reg node428_l;
    reg node429_r;
    reg node429_l;
    reg node430;
    reg node431;
    reg node432_r;
    reg node432_l;
    reg node433;
    reg node434;
    reg node435_r;
    reg node435_l;
    reg node436_r;
    reg node436_l;
    reg node437_r;
    reg node437_l;
    reg node438_r;
    reg node438_l;
    reg node439;
    reg node440;
    reg node441_r;
    reg node441_l;
    reg node442;
    reg node443;
    reg node444_r;
    reg node444_l;
    reg node445;
    reg node446;
    reg node447_r;
    reg node447_l;
    reg node448_r;
    reg node448_l;
    reg node449_r;
    reg node449_l;
    reg node450;
    reg node451;
    reg node452_r;
    reg node452_l;
    reg node453;
    reg node454;
    reg node455;
    reg node456_r;
    reg node456_l;
    reg node457_r;
    reg node457_l;
    reg node458_r;
    reg node458_l;
    reg node459_r;
    reg node459_l;
    reg node460_r;
    reg node460_l;
    reg node461;
    reg node462_r;
    reg node462_l;
    reg node463;
    reg node464;
    reg node465_r;
    reg node465_l;
    reg node466_r;
    reg node466_l;
    reg node467;
    reg node468;
    reg node469;
    reg node470_r;
    reg node470_l;
    reg node471_r;
    reg node471_l;
    reg node472_r;
    reg node472_l;
    reg node473;
    reg node474;
    reg node475_r;
    reg node475_l;
    reg node476;
    reg node477;
    reg node478_r;
    reg node478_l;
    reg node479_r;
    reg node479_l;
    reg node480;
    reg node481;
    reg node482_r;
    reg node482_l;
    reg node483;
    reg node484;
    reg node485_r;
    reg node485_l;
    reg node486_r;
    reg node486_l;
    reg node487;
    reg node488;
    reg node489_r;
    reg node489_l;
    reg node490;
    reg node491;
    reg node492_r;
    reg node492_l;
    reg node493_r;
    reg node493_l;
    reg node494_r;
    reg node494_l;
    reg node495_r;
    reg node495_l;
    reg node496_r;
    reg node496_l;
    reg node497;
    reg node498;
    reg node499_r;
    reg node499_l;
    reg node500;
    reg node501;
    reg node502_r;
    reg node502_l;
    reg node503_r;
    reg node503_l;
    reg node504;
    reg node505;
    reg node506_r;
    reg node506_l;
    reg node507;
    reg node508;
    reg node509_r;
    reg node509_l;
    reg node510;
    reg node511_r;
    reg node511_l;
    reg node512_r;
    reg node512_l;
    reg node513;
    reg node514;
    reg node515;
    reg node516_r;
    reg node516_l;
    reg node517_r;
    reg node517_l;
    reg node518_r;
    reg node518_l;
    reg node519_r;
    reg node519_l;
    reg node520;
    reg node521;
    reg node522_r;
    reg node522_l;
    reg node523;
    reg node524;
    reg node525_r;
    reg node525_l;
    reg node526_r;
    reg node526_l;
    reg node527;
    reg node528;
    reg node529;
    reg node530_r;
    reg node530_l;
    reg node531_r;
    reg node531_l;
    reg node532_r;
    reg node532_l;
    reg node533;
    reg node534;
    reg node535_r;
    reg node535_l;
    reg node536;
    reg node537;
    reg node538_r;
    reg node538_l;
    reg node539_r;
    reg node539_l;
    reg node540;
    reg node541;
    reg node542_r;
    reg node542_l;
    reg node543;
    reg node544;
    reg node545_r;
    reg node545_l;
    reg node546_r;
    reg node546_l;
    reg node547_r;
    reg node547_l;
    reg node548_r;
    reg node548_l;
    reg node549_r;
    reg node549_l;
    reg node550_r;
    reg node550_l;
    reg node551_r;
    reg node551_l;
    reg node552;
    reg node553;
    reg node554_r;
    reg node554_l;
    reg node555;
    reg node556;
    reg node557_r;
    reg node557_l;
    reg node558_r;
    reg node558_l;
    reg node559;
    reg node560;
    reg node561;
    reg node562_r;
    reg node562_l;
    reg node563;
    reg node564;
    reg node565_r;
    reg node565_l;
    reg node566_r;
    reg node566_l;
    reg node567_r;
    reg node567_l;
    reg node568_r;
    reg node568_l;
    reg node569;
    reg node570;
    reg node571_r;
    reg node571_l;
    reg node572;
    reg node573;
    reg node574_r;
    reg node574_l;
    reg node575;
    reg node576_r;
    reg node576_l;
    reg node577;
    reg node578;
    reg node579_r;
    reg node579_l;
    reg node580_r;
    reg node580_l;
    reg node581_r;
    reg node581_l;
    reg node582;
    reg node583;
    reg node584_r;
    reg node584_l;
    reg node585;
    reg node586;
    reg node587_r;
    reg node587_l;
    reg node588_r;
    reg node588_l;
    reg node589;
    reg node590;
    reg node591_r;
    reg node591_l;
    reg node592;
    reg node593;
    reg node594_r;
    reg node594_l;
    reg node595_r;
    reg node595_l;
    reg node596_r;
    reg node596_l;
    reg node597_r;
    reg node597_l;
    reg node598_r;
    reg node598_l;
    reg node599;
    reg node600;
    reg node601_r;
    reg node601_l;
    reg node602;
    reg node603;
    reg node604_r;
    reg node604_l;
    reg node605_r;
    reg node605_l;
    reg node606;
    reg node607;
    reg node608_r;
    reg node608_l;
    reg node609;
    reg node610;
    reg node611_r;
    reg node611_l;
    reg node612_r;
    reg node612_l;
    reg node613_r;
    reg node613_l;
    reg node614;
    reg node615;
    reg node616_r;
    reg node616_l;
    reg node617;
    reg node618;
    reg node619_r;
    reg node619_l;
    reg node620_r;
    reg node620_l;
    reg node621;
    reg node622;
    reg node623_r;
    reg node623_l;
    reg node624;
    reg node625;
    reg node626_r;
    reg node626_l;
    reg node627_r;
    reg node627_l;
    reg node628_r;
    reg node628_l;
    reg node629_r;
    reg node629_l;
    reg node630;
    reg node631;
    reg node632_r;
    reg node632_l;
    reg node633;
    reg node634;
    reg node635_r;
    reg node635_l;
    reg node636_r;
    reg node636_l;
    reg node637;
    reg node638;
    reg node639_r;
    reg node639_l;
    reg node640;
    reg node641;
    reg node642_r;
    reg node642_l;
    reg node643_r;
    reg node643_l;
    reg node644_r;
    reg node644_l;
    reg node645;
    reg node646;
    reg node647_r;
    reg node647_l;
    reg node648;
    reg node649;
    reg node650_r;
    reg node650_l;
    reg node651_r;
    reg node651_l;
    reg node652;
    reg node653;
    reg node654_r;
    reg node654_l;
    reg node655;
    reg node656;
    reg node657_r;
    reg node657_l;
    reg node658_r;
    reg node658_l;
    reg node659_r;
    reg node659_l;
    reg node660_r;
    reg node660_l;
    reg node661_r;
    reg node661_l;
    reg node662;
    reg node663;
    reg node664_r;
    reg node664_l;
    reg node665_r;
    reg node665_l;
    reg node666;
    reg node667;
    reg node668;
    reg node669_r;
    reg node669_l;
    reg node670_r;
    reg node670_l;
    reg node671;
    reg node672;
    reg node673_r;
    reg node673_l;
    reg node674_r;
    reg node674_l;
    reg node675;
    reg node676;
    reg node677;
    reg node678_r;
    reg node678_l;
    reg node679_r;
    reg node679_l;
    reg node680_r;
    reg node680_l;
    reg node681_r;
    reg node681_l;
    reg node682;
    reg node683;
    reg node684_r;
    reg node684_l;
    reg node685;
    reg node686;
    reg node687_r;
    reg node687_l;
    reg node688;
    reg node689;
    reg node690_r;
    reg node690_l;
    reg node691;
    reg node692_r;
    reg node692_l;
    reg node693;
    reg node694;
    reg node695_r;
    reg node695_l;
    reg node696_r;
    reg node696_l;
    reg node697_r;
    reg node697_l;
    reg node698_r;
    reg node698_l;
    reg node699_r;
    reg node699_l;
    reg node700;
    reg node701;
    reg node702;
    reg node703_r;
    reg node703_l;
    reg node704_r;
    reg node704_l;
    reg node705;
    reg node706;
    reg node707_r;
    reg node707_l;
    reg node708;
    reg node709;
    reg node710_r;
    reg node710_l;
    reg node711;
    reg node712_r;
    reg node712_l;
    reg node713;
    reg node714_r;
    reg node714_l;
    reg node715;
    reg node716;
    reg node717_r;
    reg node717_l;
    reg node718_r;
    reg node718_l;
    reg node719_r;
    reg node719_l;
    reg node720_r;
    reg node720_l;
    reg node721;
    reg node722;
    reg node723_r;
    reg node723_l;
    reg node724;
    reg node725;
    reg node726;
    reg node727_r;
    reg node727_l;
    reg node728;
    reg node729;
    reg node730_r;
    reg node730_l;
    reg node731_r;
    reg node731_l;
    reg node732_r;
    reg node732_l;
    reg node733_r;
    reg node733_l;
    reg node734_r;
    reg node734_l;
    reg node735_r;
    reg node735_l;
    reg node736_r;
    reg node736_l;
    reg node737_r;
    reg node737_l;
    reg node738_r;
    reg node738_l;
    reg node739;
    reg node740;
    reg node741_r;
    reg node741_l;
    reg node742;
    reg node743;
    reg node744_r;
    reg node744_l;
    reg node745_r;
    reg node745_l;
    reg node746;
    reg node747;
    reg node748_r;
    reg node748_l;
    reg node749;
    reg node750;
    reg node751_r;
    reg node751_l;
    reg node752_r;
    reg node752_l;
    reg node753_r;
    reg node753_l;
    reg node754;
    reg node755;
    reg node756_r;
    reg node756_l;
    reg node757;
    reg node758;
    reg node759_r;
    reg node759_l;
    reg node760_r;
    reg node760_l;
    reg node761;
    reg node762;
    reg node763_r;
    reg node763_l;
    reg node764;
    reg node765;
    reg node766_r;
    reg node766_l;
    reg node767_r;
    reg node767_l;
    reg node768_r;
    reg node768_l;
    reg node769_r;
    reg node769_l;
    reg node770;
    reg node771;
    reg node772_r;
    reg node772_l;
    reg node773;
    reg node774;
    reg node775_r;
    reg node775_l;
    reg node776_r;
    reg node776_l;
    reg node777;
    reg node778;
    reg node779_r;
    reg node779_l;
    reg node780;
    reg node781;
    reg node782_r;
    reg node782_l;
    reg node783_r;
    reg node783_l;
    reg node784_r;
    reg node784_l;
    reg node785;
    reg node786;
    reg node787_r;
    reg node787_l;
    reg node788;
    reg node789;
    reg node790_r;
    reg node790_l;
    reg node791_r;
    reg node791_l;
    reg node792;
    reg node793;
    reg node794_r;
    reg node794_l;
    reg node795;
    reg node796;
    reg node797_r;
    reg node797_l;
    reg node798_r;
    reg node798_l;
    reg node799_r;
    reg node799_l;
    reg node800_r;
    reg node800_l;
    reg node801_r;
    reg node801_l;
    reg node802;
    reg node803;
    reg node804_r;
    reg node804_l;
    reg node805;
    reg node806;
    reg node807_r;
    reg node807_l;
    reg node808_r;
    reg node808_l;
    reg node809;
    reg node810;
    reg node811_r;
    reg node811_l;
    reg node812;
    reg node813;
    reg node814_r;
    reg node814_l;
    reg node815_r;
    reg node815_l;
    reg node816_r;
    reg node816_l;
    reg node817;
    reg node818;
    reg node819_r;
    reg node819_l;
    reg node820;
    reg node821;
    reg node822;
    reg node823_r;
    reg node823_l;
    reg node824_r;
    reg node824_l;
    reg node825_r;
    reg node825_l;
    reg node826;
    reg node827_r;
    reg node827_l;
    reg node828;
    reg node829;
    reg node830_r;
    reg node830_l;
    reg node831_r;
    reg node831_l;
    reg node832;
    reg node833;
    reg node834_r;
    reg node834_l;
    reg node835;
    reg node836;
    reg node837_r;
    reg node837_l;
    reg node838_r;
    reg node838_l;
    reg node839;
    reg node840_r;
    reg node840_l;
    reg node841;
    reg node842;
    reg node843_r;
    reg node843_l;
    reg node844_r;
    reg node844_l;
    reg node845;
    reg node846;
    reg node847_r;
    reg node847_l;
    reg node848;
    reg node849;
    reg node850_r;
    reg node850_l;
    reg node851_r;
    reg node851_l;
    reg node852_r;
    reg node852_l;
    reg node853_r;
    reg node853_l;
    reg node854_r;
    reg node854_l;
    reg node855_r;
    reg node855_l;
    reg node856;
    reg node857;
    reg node858_r;
    reg node858_l;
    reg node859;
    reg node860;
    reg node861_r;
    reg node861_l;
    reg node862_r;
    reg node862_l;
    reg node863;
    reg node864;
    reg node865_r;
    reg node865_l;
    reg node866;
    reg node867;
    reg node868_r;
    reg node868_l;
    reg node869_r;
    reg node869_l;
    reg node870;
    reg node871_r;
    reg node871_l;
    reg node872;
    reg node873;
    reg node874_r;
    reg node874_l;
    reg node875_r;
    reg node875_l;
    reg node876;
    reg node877;
    reg node878_r;
    reg node878_l;
    reg node879;
    reg node880;
    reg node881_r;
    reg node881_l;
    reg node882_r;
    reg node882_l;
    reg node883_r;
    reg node883_l;
    reg node884_r;
    reg node884_l;
    reg node885;
    reg node886;
    reg node887_r;
    reg node887_l;
    reg node888;
    reg node889;
    reg node890_r;
    reg node890_l;
    reg node891_r;
    reg node891_l;
    reg node892;
    reg node893;
    reg node894_r;
    reg node894_l;
    reg node895;
    reg node896;
    reg node897_r;
    reg node897_l;
    reg node898_r;
    reg node898_l;
    reg node899_r;
    reg node899_l;
    reg node900;
    reg node901;
    reg node902;
    reg node903_r;
    reg node903_l;
    reg node904_r;
    reg node904_l;
    reg node905;
    reg node906;
    reg node907_r;
    reg node907_l;
    reg node908;
    reg node909;
    reg node910_r;
    reg node910_l;
    reg node911_r;
    reg node911_l;
    reg node912_r;
    reg node912_l;
    reg node913_r;
    reg node913_l;
    reg node914_r;
    reg node914_l;
    reg node915;
    reg node916;
    reg node917_r;
    reg node917_l;
    reg node918;
    reg node919;
    reg node920_r;
    reg node920_l;
    reg node921_r;
    reg node921_l;
    reg node922;
    reg node923;
    reg node924_r;
    reg node924_l;
    reg node925;
    reg node926;
    reg node927_r;
    reg node927_l;
    reg node928_r;
    reg node928_l;
    reg node929_r;
    reg node929_l;
    reg node930;
    reg node931;
    reg node932_r;
    reg node932_l;
    reg node933;
    reg node934;
    reg node935_r;
    reg node935_l;
    reg node936_r;
    reg node936_l;
    reg node937;
    reg node938;
    reg node939;
    reg node940_r;
    reg node940_l;
    reg node941_r;
    reg node941_l;
    reg node942_r;
    reg node942_l;
    reg node943_r;
    reg node943_l;
    reg node944;
    reg node945;
    reg node946_r;
    reg node946_l;
    reg node947;
    reg node948;
    reg node949_r;
    reg node949_l;
    reg node950;
    reg node951_r;
    reg node951_l;
    reg node952;
    reg node953;
    reg node954_r;
    reg node954_l;
    reg node955_r;
    reg node955_l;
    reg node956;
    reg node957_r;
    reg node957_l;
    reg node958;
    reg node959;
    reg node960;
    reg node961_r;
    reg node961_l;
    reg node962_r;
    reg node962_l;
    reg node963_r;
    reg node963_l;
    reg node964_r;
    reg node964_l;
    reg node965_r;
    reg node965_l;
    reg node966_r;
    reg node966_l;
    reg node967_r;
    reg node967_l;
    reg node968;
    reg node969;
    reg node970_r;
    reg node970_l;
    reg node971;
    reg node972;
    reg node973_r;
    reg node973_l;
    reg node974_r;
    reg node974_l;
    reg node975;
    reg node976;
    reg node977_r;
    reg node977_l;
    reg node978;
    reg node979;
    reg node980_r;
    reg node980_l;
    reg node981_r;
    reg node981_l;
    reg node982_r;
    reg node982_l;
    reg node983;
    reg node984;
    reg node985_r;
    reg node985_l;
    reg node986;
    reg node987;
    reg node988_r;
    reg node988_l;
    reg node989_r;
    reg node989_l;
    reg node990;
    reg node991;
    reg node992_r;
    reg node992_l;
    reg node993;
    reg node994;
    reg node995_r;
    reg node995_l;
    reg node996_r;
    reg node996_l;
    reg node997_r;
    reg node997_l;
    reg node998_r;
    reg node998_l;
    reg node999;
    reg node1000;
    reg node1001_r;
    reg node1001_l;
    reg node1002;
    reg node1003;
    reg node1004_r;
    reg node1004_l;
    reg node1005;
    reg node1006;
    reg node1007_r;
    reg node1007_l;
    reg node1008_r;
    reg node1008_l;
    reg node1009;
    reg node1010_r;
    reg node1010_l;
    reg node1011;
    reg node1012;
    reg node1013_r;
    reg node1013_l;
    reg node1014_r;
    reg node1014_l;
    reg node1015;
    reg node1016;
    reg node1017_r;
    reg node1017_l;
    reg node1018;
    reg node1019;
    reg node1020_r;
    reg node1020_l;
    reg node1021_r;
    reg node1021_l;
    reg node1022_r;
    reg node1022_l;
    reg node1023_r;
    reg node1023_l;
    reg node1024_r;
    reg node1024_l;
    reg node1025;
    reg node1026;
    reg node1027_r;
    reg node1027_l;
    reg node1028;
    reg node1029;
    reg node1030_r;
    reg node1030_l;
    reg node1031_r;
    reg node1031_l;
    reg node1032;
    reg node1033;
    reg node1034_r;
    reg node1034_l;
    reg node1035;
    reg node1036;
    reg node1037_r;
    reg node1037_l;
    reg node1038_r;
    reg node1038_l;
    reg node1039_r;
    reg node1039_l;
    reg node1040;
    reg node1041;
    reg node1042_r;
    reg node1042_l;
    reg node1043;
    reg node1044;
    reg node1045_r;
    reg node1045_l;
    reg node1046_r;
    reg node1046_l;
    reg node1047;
    reg node1048;
    reg node1049_r;
    reg node1049_l;
    reg node1050;
    reg node1051;
    reg node1052_r;
    reg node1052_l;
    reg node1053_r;
    reg node1053_l;
    reg node1054_r;
    reg node1054_l;
    reg node1055_r;
    reg node1055_l;
    reg node1056;
    reg node1057;
    reg node1058_r;
    reg node1058_l;
    reg node1059;
    reg node1060;
    reg node1061_r;
    reg node1061_l;
    reg node1062_r;
    reg node1062_l;
    reg node1063;
    reg node1064;
    reg node1065_r;
    reg node1065_l;
    reg node1066;
    reg node1067;
    reg node1068_r;
    reg node1068_l;
    reg node1069_r;
    reg node1069_l;
    reg node1070_r;
    reg node1070_l;
    reg node1071;
    reg node1072;
    reg node1073_r;
    reg node1073_l;
    reg node1074;
    reg node1075;
    reg node1076_r;
    reg node1076_l;
    reg node1077_r;
    reg node1077_l;
    reg node1078;
    reg node1079;
    reg node1080_r;
    reg node1080_l;
    reg node1081;
    reg node1082;
    reg node1083_r;
    reg node1083_l;
    reg node1084_r;
    reg node1084_l;
    reg node1085_r;
    reg node1085_l;
    reg node1086_r;
    reg node1086_l;
    reg node1087_r;
    reg node1087_l;
    reg node1088_r;
    reg node1088_l;
    reg node1089;
    reg node1090;
    reg node1091_r;
    reg node1091_l;
    reg node1092;
    reg node1093;
    reg node1094_r;
    reg node1094_l;
    reg node1095_r;
    reg node1095_l;
    reg node1096;
    reg node1097;
    reg node1098_r;
    reg node1098_l;
    reg node1099;
    reg node1100;
    reg node1101_r;
    reg node1101_l;
    reg node1102_r;
    reg node1102_l;
    reg node1103_r;
    reg node1103_l;
    reg node1104;
    reg node1105;
    reg node1106;
    reg node1107_r;
    reg node1107_l;
    reg node1108_r;
    reg node1108_l;
    reg node1109;
    reg node1110;
    reg node1111_r;
    reg node1111_l;
    reg node1112;
    reg node1113;
    reg node1114_r;
    reg node1114_l;
    reg node1115_r;
    reg node1115_l;
    reg node1116_r;
    reg node1116_l;
    reg node1117_r;
    reg node1117_l;
    reg node1118;
    reg node1119;
    reg node1120_r;
    reg node1120_l;
    reg node1121;
    reg node1122;
    reg node1123_r;
    reg node1123_l;
    reg node1124;
    reg node1125_r;
    reg node1125_l;
    reg node1126;
    reg node1127;
    reg node1128_r;
    reg node1128_l;
    reg node1129_r;
    reg node1129_l;
    reg node1130_r;
    reg node1130_l;
    reg node1131;
    reg node1132;
    reg node1133;
    reg node1134_r;
    reg node1134_l;
    reg node1135_r;
    reg node1135_l;
    reg node1136;
    reg node1137;
    reg node1138;
    reg node1139_r;
    reg node1139_l;
    reg node1140_r;
    reg node1140_l;
    reg node1141_r;
    reg node1141_l;
    reg node1142_r;
    reg node1142_l;
    reg node1143_r;
    reg node1143_l;
    reg node1144;
    reg node1145;
    reg node1146_r;
    reg node1146_l;
    reg node1147;
    reg node1148;
    reg node1149_r;
    reg node1149_l;
    reg node1150_r;
    reg node1150_l;
    reg node1151;
    reg node1152;
    reg node1153_r;
    reg node1153_l;
    reg node1154;
    reg node1155;
    reg node1156_r;
    reg node1156_l;
    reg node1157_r;
    reg node1157_l;
    reg node1158_r;
    reg node1158_l;
    reg node1159;
    reg node1160;
    reg node1161_r;
    reg node1161_l;
    reg node1162;
    reg node1163;
    reg node1164_r;
    reg node1164_l;
    reg node1165_r;
    reg node1165_l;
    reg node1166;
    reg node1167;
    reg node1168_r;
    reg node1168_l;
    reg node1169;
    reg node1170;
    reg node1171_r;
    reg node1171_l;
    reg node1172_r;
    reg node1172_l;
    reg node1173_r;
    reg node1173_l;
    reg node1174_r;
    reg node1174_l;
    reg node1175;
    reg node1176;
    reg node1177;
    reg node1178_r;
    reg node1178_l;
    reg node1179_r;
    reg node1179_l;
    reg node1180;
    reg node1181;
    reg node1182_r;
    reg node1182_l;
    reg node1183;
    reg node1184;
    reg node1185_r;
    reg node1185_l;
    reg node1186_r;
    reg node1186_l;
    reg node1187_r;
    reg node1187_l;
    reg node1188;
    reg node1189;
    reg node1190_r;
    reg node1190_l;
    reg node1191;
    reg node1192;
    reg node1193_r;
    reg node1193_l;
    reg node1194_r;
    reg node1194_l;
    reg node1195;
    reg node1196;
    reg node1197_r;
    reg node1197_l;
    reg node1198;
    reg node1199;
    reg node1200_r;
    reg node1200_l;
    reg node1201_r;
    reg node1201_l;
    reg node1202_r;
    reg node1202_l;
    reg node1203_r;
    reg node1203_l;
    reg node1204_r;
    reg node1204_l;
    reg node1205_r;
    reg node1205_l;
    reg node1206_r;
    reg node1206_l;
    reg node1207_r;
    reg node1207_l;
    reg node1208;
    reg node1209;
    reg node1210_r;
    reg node1210_l;
    reg node1211;
    reg node1212;
    reg node1213_r;
    reg node1213_l;
    reg node1214_r;
    reg node1214_l;
    reg node1215;
    reg node1216;
    reg node1217_r;
    reg node1217_l;
    reg node1218;
    reg node1219;
    reg node1220_r;
    reg node1220_l;
    reg node1221_r;
    reg node1221_l;
    reg node1222_r;
    reg node1222_l;
    reg node1223;
    reg node1224;
    reg node1225_r;
    reg node1225_l;
    reg node1226;
    reg node1227;
    reg node1228_r;
    reg node1228_l;
    reg node1229_r;
    reg node1229_l;
    reg node1230;
    reg node1231;
    reg node1232_r;
    reg node1232_l;
    reg node1233;
    reg node1234;
    reg node1235_r;
    reg node1235_l;
    reg node1236_r;
    reg node1236_l;
    reg node1237_r;
    reg node1237_l;
    reg node1238_r;
    reg node1238_l;
    reg node1239;
    reg node1240;
    reg node1241_r;
    reg node1241_l;
    reg node1242;
    reg node1243;
    reg node1244_r;
    reg node1244_l;
    reg node1245_r;
    reg node1245_l;
    reg node1246;
    reg node1247;
    reg node1248_r;
    reg node1248_l;
    reg node1249;
    reg node1250;
    reg node1251_r;
    reg node1251_l;
    reg node1252_r;
    reg node1252_l;
    reg node1253_r;
    reg node1253_l;
    reg node1254;
    reg node1255;
    reg node1256_r;
    reg node1256_l;
    reg node1257;
    reg node1258;
    reg node1259_r;
    reg node1259_l;
    reg node1260_r;
    reg node1260_l;
    reg node1261;
    reg node1262;
    reg node1263_r;
    reg node1263_l;
    reg node1264;
    reg node1265;
    reg node1266_r;
    reg node1266_l;
    reg node1267_r;
    reg node1267_l;
    reg node1268_r;
    reg node1268_l;
    reg node1269_r;
    reg node1269_l;
    reg node1270_r;
    reg node1270_l;
    reg node1271;
    reg node1272;
    reg node1273;
    reg node1274_r;
    reg node1274_l;
    reg node1275_r;
    reg node1275_l;
    reg node1276;
    reg node1277;
    reg node1278_r;
    reg node1278_l;
    reg node1279;
    reg node1280;
    reg node1281_r;
    reg node1281_l;
    reg node1282_r;
    reg node1282_l;
    reg node1283_r;
    reg node1283_l;
    reg node1284;
    reg node1285;
    reg node1286_r;
    reg node1286_l;
    reg node1287;
    reg node1288;
    reg node1289_r;
    reg node1289_l;
    reg node1290_r;
    reg node1290_l;
    reg node1291;
    reg node1292;
    reg node1293_r;
    reg node1293_l;
    reg node1294;
    reg node1295;
    reg node1296_r;
    reg node1296_l;
    reg node1297_r;
    reg node1297_l;
    reg node1298_r;
    reg node1298_l;
    reg node1299_r;
    reg node1299_l;
    reg node1300;
    reg node1301;
    reg node1302_r;
    reg node1302_l;
    reg node1303;
    reg node1304;
    reg node1305_r;
    reg node1305_l;
    reg node1306_r;
    reg node1306_l;
    reg node1307;
    reg node1308;
    reg node1309;
    reg node1310_r;
    reg node1310_l;
    reg node1311_r;
    reg node1311_l;
    reg node1312_r;
    reg node1312_l;
    reg node1313;
    reg node1314;
    reg node1315_r;
    reg node1315_l;
    reg node1316;
    reg node1317;
    reg node1318_r;
    reg node1318_l;
    reg node1319;
    reg node1320;
    reg node1321_r;
    reg node1321_l;
    reg node1322_r;
    reg node1322_l;
    reg node1323_r;
    reg node1323_l;
    reg node1324_r;
    reg node1324_l;
    reg node1325_r;
    reg node1325_l;
    reg node1326_r;
    reg node1326_l;
    reg node1327;
    reg node1328;
    reg node1329_r;
    reg node1329_l;
    reg node1330;
    reg node1331;
    reg node1332_r;
    reg node1332_l;
    reg node1333_r;
    reg node1333_l;
    reg node1334;
    reg node1335;
    reg node1336_r;
    reg node1336_l;
    reg node1337;
    reg node1338;
    reg node1339_r;
    reg node1339_l;
    reg node1340_r;
    reg node1340_l;
    reg node1341_r;
    reg node1341_l;
    reg node1342;
    reg node1343;
    reg node1344_r;
    reg node1344_l;
    reg node1345;
    reg node1346;
    reg node1347_r;
    reg node1347_l;
    reg node1348_r;
    reg node1348_l;
    reg node1349;
    reg node1350;
    reg node1351_r;
    reg node1351_l;
    reg node1352;
    reg node1353;
    reg node1354_r;
    reg node1354_l;
    reg node1355_r;
    reg node1355_l;
    reg node1356;
    reg node1357_r;
    reg node1357_l;
    reg node1358_r;
    reg node1358_l;
    reg node1359;
    reg node1360;
    reg node1361;
    reg node1362_r;
    reg node1362_l;
    reg node1363_r;
    reg node1363_l;
    reg node1364_r;
    reg node1364_l;
    reg node1365;
    reg node1366;
    reg node1367_r;
    reg node1367_l;
    reg node1368;
    reg node1369;
    reg node1370_r;
    reg node1370_l;
    reg node1371;
    reg node1372;
    reg node1373_r;
    reg node1373_l;
    reg node1374_r;
    reg node1374_l;
    reg node1375_r;
    reg node1375_l;
    reg node1376_r;
    reg node1376_l;
    reg node1377;
    reg node1378_r;
    reg node1378_l;
    reg node1379;
    reg node1380;
    reg node1381_r;
    reg node1381_l;
    reg node1382_r;
    reg node1382_l;
    reg node1383;
    reg node1384;
    reg node1385_r;
    reg node1385_l;
    reg node1386;
    reg node1387;
    reg node1388_r;
    reg node1388_l;
    reg node1389_r;
    reg node1389_l;
    reg node1390;
    reg node1391;
    reg node1392_r;
    reg node1392_l;
    reg node1393_r;
    reg node1393_l;
    reg node1394;
    reg node1395;
    reg node1396;
    reg node1397_r;
    reg node1397_l;
    reg node1398_r;
    reg node1398_l;
    reg node1399;
    reg node1400_r;
    reg node1400_l;
    reg node1401_r;
    reg node1401_l;
    reg node1402;
    reg node1403;
    reg node1404_r;
    reg node1404_l;
    reg node1405;
    reg node1406;
    reg node1407_r;
    reg node1407_l;
    reg node1408_r;
    reg node1408_l;
    reg node1409;
    reg node1410;
    reg node1411_r;
    reg node1411_l;
    reg node1412_r;
    reg node1412_l;
    reg node1413;
    reg node1414;
    reg node1415;
    reg node1416_r;
    reg node1416_l;
    reg node1417_r;
    reg node1417_l;
    reg node1418_r;
    reg node1418_l;
    reg node1419_r;
    reg node1419_l;
    reg node1420_r;
    reg node1420_l;
    reg node1421_r;
    reg node1421_l;
    reg node1422_r;
    reg node1422_l;
    reg node1423;
    reg node1424;
    reg node1425_r;
    reg node1425_l;
    reg node1426;
    reg node1427;
    reg node1428_r;
    reg node1428_l;
    reg node1429_r;
    reg node1429_l;
    reg node1430;
    reg node1431;
    reg node1432_r;
    reg node1432_l;
    reg node1433;
    reg node1434;
    reg node1435_r;
    reg node1435_l;
    reg node1436_r;
    reg node1436_l;
    reg node1437_r;
    reg node1437_l;
    reg node1438;
    reg node1439;
    reg node1440_r;
    reg node1440_l;
    reg node1441;
    reg node1442;
    reg node1443_r;
    reg node1443_l;
    reg node1444;
    reg node1445_r;
    reg node1445_l;
    reg node1446;
    reg node1447;
    reg node1448_r;
    reg node1448_l;
    reg node1449_r;
    reg node1449_l;
    reg node1450_r;
    reg node1450_l;
    reg node1451_r;
    reg node1451_l;
    reg node1452;
    reg node1453;
    reg node1454_r;
    reg node1454_l;
    reg node1455;
    reg node1456;
    reg node1457_r;
    reg node1457_l;
    reg node1458_r;
    reg node1458_l;
    reg node1459;
    reg node1460;
    reg node1461_r;
    reg node1461_l;
    reg node1462;
    reg node1463;
    reg node1464_r;
    reg node1464_l;
    reg node1465_r;
    reg node1465_l;
    reg node1466_r;
    reg node1466_l;
    reg node1467;
    reg node1468;
    reg node1469_r;
    reg node1469_l;
    reg node1470;
    reg node1471;
    reg node1472_r;
    reg node1472_l;
    reg node1473_r;
    reg node1473_l;
    reg node1474;
    reg node1475;
    reg node1476_r;
    reg node1476_l;
    reg node1477;
    reg node1478;
    reg node1479_r;
    reg node1479_l;
    reg node1480_r;
    reg node1480_l;
    reg node1481_r;
    reg node1481_l;
    reg node1482_r;
    reg node1482_l;
    reg node1483_r;
    reg node1483_l;
    reg node1484;
    reg node1485;
    reg node1486_r;
    reg node1486_l;
    reg node1487;
    reg node1488;
    reg node1489_r;
    reg node1489_l;
    reg node1490_r;
    reg node1490_l;
    reg node1491;
    reg node1492;
    reg node1493_r;
    reg node1493_l;
    reg node1494;
    reg node1495;
    reg node1496_r;
    reg node1496_l;
    reg node1497_r;
    reg node1497_l;
    reg node1498;
    reg node1499_r;
    reg node1499_l;
    reg node1500;
    reg node1501;
    reg node1502_r;
    reg node1502_l;
    reg node1503_r;
    reg node1503_l;
    reg node1504;
    reg node1505;
    reg node1506;
    reg node1507_r;
    reg node1507_l;
    reg node1508_r;
    reg node1508_l;
    reg node1509;
    reg node1510_r;
    reg node1510_l;
    reg node1511_r;
    reg node1511_l;
    reg node1512;
    reg node1513;
    reg node1514_r;
    reg node1514_l;
    reg node1515;
    reg node1516;
    reg node1517_r;
    reg node1517_l;
    reg node1518_r;
    reg node1518_l;
    reg node1519_r;
    reg node1519_l;
    reg node1520;
    reg node1521;
    reg node1522_r;
    reg node1522_l;
    reg node1523;
    reg node1524;
    reg node1525_r;
    reg node1525_l;
    reg node1526_r;
    reg node1526_l;
    reg node1527;
    reg node1528;
    reg node1529_r;
    reg node1529_l;
    reg node1530;
    reg node1531;
    reg node1532_r;
    reg node1532_l;
    reg node1533_r;
    reg node1533_l;
    reg node1534_r;
    reg node1534_l;
    reg node1535_r;
    reg node1535_l;
    reg node1536_r;
    reg node1536_l;
    reg node1537_r;
    reg node1537_l;
    reg node1538;
    reg node1539;
    reg node1540_r;
    reg node1540_l;
    reg node1541;
    reg node1542;
    reg node1543_r;
    reg node1543_l;
    reg node1544_r;
    reg node1544_l;
    reg node1545;
    reg node1546;
    reg node1547_r;
    reg node1547_l;
    reg node1548;
    reg node1549;
    reg node1550_r;
    reg node1550_l;
    reg node1551_r;
    reg node1551_l;
    reg node1552_r;
    reg node1552_l;
    reg node1553;
    reg node1554;
    reg node1555_r;
    reg node1555_l;
    reg node1556;
    reg node1557;
    reg node1558_r;
    reg node1558_l;
    reg node1559_r;
    reg node1559_l;
    reg node1560;
    reg node1561;
    reg node1562;
    reg node1563_r;
    reg node1563_l;
    reg node1564_r;
    reg node1564_l;
    reg node1565_r;
    reg node1565_l;
    reg node1566_r;
    reg node1566_l;
    reg node1567;
    reg node1568;
    reg node1569_r;
    reg node1569_l;
    reg node1570;
    reg node1571;
    reg node1572_r;
    reg node1572_l;
    reg node1573_r;
    reg node1573_l;
    reg node1574;
    reg node1575;
    reg node1576_r;
    reg node1576_l;
    reg node1577;
    reg node1578;
    reg node1579_r;
    reg node1579_l;
    reg node1580_r;
    reg node1580_l;
    reg node1581_r;
    reg node1581_l;
    reg node1582;
    reg node1583;
    reg node1584_r;
    reg node1584_l;
    reg node1585;
    reg node1586;
    reg node1587_r;
    reg node1587_l;
    reg node1588_r;
    reg node1588_l;
    reg node1589;
    reg node1590;
    reg node1591;
    reg node1592_r;
    reg node1592_l;
    reg node1593_r;
    reg node1593_l;
    reg node1594_r;
    reg node1594_l;
    reg node1595_r;
    reg node1595_l;
    reg node1596_r;
    reg node1596_l;
    reg node1597;
    reg node1598;
    reg node1599_r;
    reg node1599_l;
    reg node1600;
    reg node1601;
    reg node1602_r;
    reg node1602_l;
    reg node1603_r;
    reg node1603_l;
    reg node1604;
    reg node1605;
    reg node1606_r;
    reg node1606_l;
    reg node1607;
    reg node1608;
    reg node1609_r;
    reg node1609_l;
    reg node1610_r;
    reg node1610_l;
    reg node1611_r;
    reg node1611_l;
    reg node1612;
    reg node1613;
    reg node1614_r;
    reg node1614_l;
    reg node1615;
    reg node1616;
    reg node1617_r;
    reg node1617_l;
    reg node1618_r;
    reg node1618_l;
    reg node1619;
    reg node1620;
    reg node1621_r;
    reg node1621_l;
    reg node1622;
    reg node1623;
    reg node1624_r;
    reg node1624_l;
    reg node1625_r;
    reg node1625_l;
    reg node1626_r;
    reg node1626_l;
    reg node1627_r;
    reg node1627_l;
    reg node1628;
    reg node1629;
    reg node1630_r;
    reg node1630_l;
    reg node1631;
    reg node1632;
    reg node1633_r;
    reg node1633_l;
    reg node1634_r;
    reg node1634_l;
    reg node1635;
    reg node1636;
    reg node1637_r;
    reg node1637_l;
    reg node1638;
    reg node1639;
    reg node1640_r;
    reg node1640_l;
    reg node1641_r;
    reg node1641_l;
    reg node1642_r;
    reg node1642_l;
    reg node1643;
    reg node1644;
    reg node1645_r;
    reg node1645_l;
    reg node1646;
    reg node1647;
    reg node1648_r;
    reg node1648_l;
    reg node1649_r;
    reg node1649_l;
    reg node1650;
    reg node1651;
    reg node1652;
    reg result0;
    reg result1;
    reg result2;
    reg result3;
    reg result4;
    reg result5;
    reg result6;
    reg result7;
    reg result8;
    reg result9;

    begin
      node0_r = pixel[378];
      node0_l = ~pixel[378];
      node1_r = node0_l & pixel[539];
      node1_l = node0_l & ~pixel[539];
      node2_r = node1_l & pixel[433];
      node2_l = node1_l & ~pixel[433];
      node3_r = node2_l & pixel[541];
      node3_l = node2_l & ~pixel[541];
      node4_r = node3_l & pixel[457];
      node4_l = node3_l & ~pixel[457];
      node5_r = node4_l & pixel[183];
      node5_l = node4_l & ~pixel[183];
      node6_r = node5_l & pixel[404];
      node6_l = node5_l & ~pixel[404];
      node7_r = node6_l & pixel[128];
      node7_l = node6_l & ~pixel[128];
      node8_r = node7_l & pixel[469];
      node8_l = node7_l & ~pixel[469];
      node9_r = node8_l & pixel[460];
      node9_l = node8_l & ~pixel[460];
      node10 = node9_l;
      node11 = node9_r;
      node12_r = node8_r & pixel[537];
      node12_l = node8_r & ~pixel[537];
      node13 = node12_l;
      node14 = node12_r;
      node15_r = node7_r & pixel[403];
      node15_l = node7_r & ~pixel[403];
      node16_r = node15_l & pixel[270];
      node16_l = node15_l & ~pixel[270];
      node17 = node16_l;
      node18 = node16_r;
      node19_r = node15_r & pixel[159];
      node19_l = node15_r & ~pixel[159];
      node20 = node19_l;
      node21 = node19_r;
      node22_r = node6_r & pixel[326];
      node22_l = node6_r & ~pixel[326];
      node23_r = node22_l & pixel[459];
      node23_l = node22_l & ~pixel[459];
      node24_r = node23_l & pixel[428];
      node24_l = node23_l & ~pixel[428];
      node25 = node24_l;
      node26 = node24_r;
      node27_r = node23_r & pixel[269];
      node27_l = node23_r & ~pixel[269];
      node28 = node27_l;
      node29 = node27_r;
      node30_r = node22_r & pixel[264];
      node30_l = node22_r & ~pixel[264];
      node31_r = node30_l & pixel[464];
      node31_l = node30_l & ~pixel[464];
      node32 = node31_l;
      node33 = node31_r;
      node34_r = node30_r & pixel[486];
      node34_l = node30_r & ~pixel[486];
      node35 = node34_l;
      node36 = node34_r;
      node37_r = node5_r & pixel[359];
      node37_l = node5_r & ~pixel[359];
      node38_r = node37_l & pixel[546];
      node38_l = node37_l & ~pixel[546];
      node39_r = node38_l & pixel[322];
      node39_l = node38_l & ~pixel[322];
      node40_r = node39_l & pixel[241];
      node40_l = node39_l & ~pixel[241];
      node41 = node40_l;
      node42 = node40_r;
      node43_r = node39_r & pixel[401];
      node43_l = node39_r & ~pixel[401];
      node44 = node43_l;
      node45 = node43_r;
      node46_r = node38_r & pixel[348];
      node46_l = node38_r & ~pixel[348];
      node47_r = node46_l & pixel[151];
      node47_l = node46_l & ~pixel[151];
      node48 = node47_l;
      node49 = node47_r;
      node50_r = node46_r & pixel[488];
      node50_l = node46_r & ~pixel[488];
      node51 = node50_l;
      node52 = node50_r;
      node53_r = node37_r & pixel[565];
      node53_l = node37_r & ~pixel[565];
      node54_r = node53_l & pixel[409];
      node54_l = node53_l & ~pixel[409];
      node55 = node54_l;
      node56 = node54_r;
      node57_r = node53_r & pixel[410];
      node57_l = node53_r & ~pixel[410];
      node58 = node57_l;
      node59_r = node57_r & pixel[524];
      node59_l = node57_r & ~pixel[524];
      node60 = node59_l;
      node61 = node59_r;
      node62_r = node4_r & pixel[99];
      node62_l = node4_r & ~pixel[99];
      node63_r = node62_l & pixel[465];
      node63_l = node62_l & ~pixel[465];
      node64_r = node63_l & pixel[413];
      node64_l = node63_l & ~pixel[413];
      node65_r = node64_l & pixel[495];
      node65_l = node64_l & ~pixel[495];
      node66_r = node65_l & pixel[380];
      node66_l = node65_l & ~pixel[380];
      node67 = node66_l;
      node68 = node66_r;
      node69_r = node65_r & pixel[487];
      node69_l = node65_r & ~pixel[487];
      node70 = node69_l;
      node71 = node69_r;
      node72_r = node64_r & pixel[518];
      node72_l = node64_r & ~pixel[518];
      node73_r = node72_l & pixel[186];
      node73_l = node72_l & ~pixel[186];
      node74 = node73_l;
      node75 = node73_r;
      node76_r = node72_r & pixel[368];
      node76_l = node72_r & ~pixel[368];
      node77 = node76_l;
      node78 = node76_r;
      node79_r = node63_r & pixel[487];
      node79_l = node63_r & ~pixel[487];
      node80_r = node79_l & pixel[152];
      node80_l = node79_l & ~pixel[152];
      node81_r = node80_l & pixel[569];
      node81_l = node80_l & ~pixel[569];
      node82 = node81_l;
      node83 = node81_r;
      node84_r = node80_r & pixel[576];
      node84_l = node80_r & ~pixel[576];
      node85 = node84_l;
      node86 = node84_r;
      node87_r = node79_r & pixel[525];
      node87_l = node79_r & ~pixel[525];
      node88_r = node87_l & pixel[183];
      node88_l = node87_l & ~pixel[183];
      node89 = node88_l;
      node90 = node88_r;
      node91_r = node87_r & pixel[665];
      node91_l = node87_r & ~pixel[665];
      node92 = node91_l;
      node93 = node91_r;
      node94_r = node62_r & pixel[264];
      node94_l = node62_r & ~pixel[264];
      node95_r = node94_l & pixel[481];
      node95_l = node94_l & ~pixel[481];
      node96_r = node95_l & pixel[214];
      node96_l = node95_l & ~pixel[214];
      node97_r = node96_l & pixel[345];
      node97_l = node96_l & ~pixel[345];
      node98 = node97_l;
      node99 = node97_r;
      node100_r = node96_r & pixel[272];
      node100_l = node96_r & ~pixel[272];
      node101 = node100_l;
      node102 = node100_r;
      node103 = node95_r;
      node104_r = node94_r & pixel[537];
      node104_l = node94_r & ~pixel[537];
      node105_r = node104_l & pixel[491];
      node105_l = node104_l & ~pixel[491];
      node106_r = node105_l & pixel[240];
      node106_l = node105_l & ~pixel[240];
      node107 = node106_l;
      node108 = node106_r;
      node109_r = node105_r & pixel[323];
      node109_l = node105_r & ~pixel[323];
      node110 = node109_l;
      node111 = node109_r;
      node112 = node104_r;
      node113_r = node3_r & pixel[516];
      node113_l = node3_r & ~pixel[516];
      node114_r = node113_l & pixel[657];
      node114_l = node113_l & ~pixel[657];
      node115_r = node114_l & pixel[627];
      node115_l = node114_l & ~pixel[627];
      node116_r = node115_l & pixel[576];
      node116_l = node115_l & ~pixel[576];
      node117_r = node116_l & pixel[329];
      node117_l = node116_l & ~pixel[329];
      node118_r = node117_l & pixel[370];
      node118_l = node117_l & ~pixel[370];
      node119 = node118_l;
      node120 = node118_r;
      node121_r = node117_r & pixel[716];
      node121_l = node117_r & ~pixel[716];
      node122 = node121_l;
      node123 = node121_r;
      node124_r = node116_r & pixel[599];
      node124_l = node116_r & ~pixel[599];
      node125_r = node124_l & pixel[573];
      node125_l = node124_l & ~pixel[573];
      node126 = node125_l;
      node127 = node125_r;
      node128_r = node124_r & pixel[268];
      node128_l = node124_r & ~pixel[268];
      node129 = node128_l;
      node130 = node128_r;
      node131_r = node115_r & pixel[435];
      node131_l = node115_r & ~pixel[435];
      node132_r = node131_l & pixel[294];
      node132_l = node131_l & ~pixel[294];
      node133_r = node132_l & pixel[607];
      node133_l = node132_l & ~pixel[607];
      node134 = node133_l;
      node135 = node133_r;
      node136_r = node132_r & pixel[318];
      node136_l = node132_r & ~pixel[318];
      node137 = node136_l;
      node138 = node136_r;
      node139_r = node131_r & pixel[603];
      node139_l = node131_r & ~pixel[603];
      node140_r = node139_l & pixel[103];
      node140_l = node139_l & ~pixel[103];
      node141 = node140_l;
      node142 = node140_r;
      node143_r = node139_r & pixel[458];
      node143_l = node139_r & ~pixel[458];
      node144 = node143_l;
      node145 = node143_r;
      node146_r = node114_r & pixel[623];
      node146_l = node114_r & ~pixel[623];
      node147_r = node146_l & pixel[349];
      node147_l = node146_l & ~pixel[349];
      node148_r = node147_l & pixel[352];
      node148_l = node147_l & ~pixel[352];
      node149_r = node148_l & pixel[570];
      node149_l = node148_l & ~pixel[570];
      node150 = node149_l;
      node151 = node149_r;
      node152_r = node148_r & pixel[457];
      node152_l = node148_r & ~pixel[457];
      node153 = node152_l;
      node154 = node152_r;
      node155_r = node147_r & pixel[178];
      node155_l = node147_r & ~pixel[178];
      node156_r = node155_l & pixel[430];
      node156_l = node155_l & ~pixel[430];
      node157 = node156_l;
      node158 = node156_r;
      node159_r = node155_r & pixel[234];
      node159_l = node155_r & ~pixel[234];
      node160 = node159_l;
      node161 = node159_r;
      node162_r = node146_r & pixel[348];
      node162_l = node146_r & ~pixel[348];
      node163 = node162_l;
      node164_r = node162_r & pixel[401];
      node164_l = node162_r & ~pixel[401];
      node165 = node164_l;
      node166_r = node164_r & pixel[270];
      node166_l = node164_r & ~pixel[270];
      node167 = node166_l;
      node168 = node166_r;
      node169_r = node113_r & pixel[102];
      node169_l = node113_r & ~pixel[102];
      node170_r = node169_l & pixel[599];
      node170_l = node169_l & ~pixel[599];
      node171_r = node170_l & pixel[240];
      node171_l = node170_l & ~pixel[240];
      node172_r = node171_l & pixel[98];
      node172_l = node171_l & ~pixel[98];
      node173_r = node172_l & pixel[442];
      node173_l = node172_l & ~pixel[442];
      node174 = node173_l;
      node175 = node173_r;
      node176_r = node172_r & pixel[468];
      node176_l = node172_r & ~pixel[468];
      node177 = node176_l;
      node178 = node176_r;
      node179_r = node171_r & pixel[327];
      node179_l = node171_r & ~pixel[327];
      node180_r = node179_l & pixel[556];
      node180_l = node179_l & ~pixel[556];
      node181 = node180_l;
      node182 = node180_r;
      node183_r = node179_r & pixel[465];
      node183_l = node179_r & ~pixel[465];
      node184 = node183_l;
      node185 = node183_r;
      node186_r = node170_r & pixel[212];
      node186_l = node170_r & ~pixel[212];
      node187_r = node186_l & pixel[654];
      node187_l = node186_l & ~pixel[654];
      node188_r = node187_l & pixel[597];
      node188_l = node187_l & ~pixel[597];
      node189 = node188_l;
      node190 = node188_r;
      node191_r = node187_r & pixel[491];
      node191_l = node187_r & ~pixel[491];
      node192 = node191_l;
      node193 = node191_r;
      node194_r = node186_r & pixel[491];
      node194_l = node186_r & ~pixel[491];
      node195_r = node194_l & pixel[571];
      node195_l = node194_l & ~pixel[571];
      node196 = node195_l;
      node197 = node195_r;
      node198_r = node194_r & pixel[580];
      node198_l = node194_r & ~pixel[580];
      node199 = node198_l;
      node200 = node198_r;
      node201_r = node169_r & pixel[298];
      node201_l = node169_r & ~pixel[298];
      node202_r = node201_l & pixel[324];
      node202_l = node201_l & ~pixel[324];
      node203_r = node202_l & pixel[301];
      node203_l = node202_l & ~pixel[301];
      node204 = node203_l;
      node205_r = node203_r & pixel[484];
      node205_l = node203_r & ~pixel[484];
      node206 = node205_l;
      node207 = node205_r;
      node208 = node202_r;
      node209_r = node201_r & pixel[348];
      node209_l = node201_r & ~pixel[348];
      node210_r = node209_l & pixel[93];
      node210_l = node209_l & ~pixel[93];
      node211 = node210_l;
      node212 = node210_r;
      node213_r = node209_r & pixel[179];
      node213_l = node209_r & ~pixel[179];
      node214_r = node213_l & pixel[576];
      node214_l = node213_l & ~pixel[576];
      node215 = node214_l;
      node216 = node214_r;
      node217 = node213_r;
      node218_r = node2_r & pixel[99];
      node218_l = node2_r & ~pixel[99];
      node219_r = node218_l & pixel[212];
      node219_l = node218_l & ~pixel[212];
      node220_r = node219_l & pixel[70];
      node220_l = node219_l & ~pixel[70];
      node221_r = node220_l & pixel[155];
      node221_l = node220_l & ~pixel[155];
      node222_r = node221_l & pixel[95];
      node222_l = node221_l & ~pixel[95];
      node223_r = node222_l & pixel[624];
      node223_l = node222_l & ~pixel[624];
      node224_r = node223_l & pixel[215];
      node224_l = node223_l & ~pixel[215];
      node225 = node224_l;
      node226 = node224_r;
      node227_r = node223_r & pixel[517];
      node227_l = node223_r & ~pixel[517];
      node228 = node227_l;
      node229 = node227_r;
      node230_r = node222_r & pixel[240];
      node230_l = node222_r & ~pixel[240];
      node231_r = node230_l & pixel[238];
      node231_l = node230_l & ~pixel[238];
      node232 = node231_l;
      node233 = node231_r;
      node234_r = node230_r & pixel[273];
      node234_l = node230_r & ~pixel[273];
      node235 = node234_l;
      node236 = node234_r;
      node237_r = node221_r & pixel[623];
      node237_l = node221_r & ~pixel[623];
      node238_r = node237_l & pixel[491];
      node238_l = node237_l & ~pixel[491];
      node239_r = node238_l & pixel[659];
      node239_l = node238_l & ~pixel[659];
      node240 = node239_l;
      node241 = node239_r;
      node242_r = node238_r & pixel[632];
      node242_l = node238_r & ~pixel[632];
      node243 = node242_l;
      node244 = node242_r;
      node245_r = node237_r & pixel[291];
      node245_l = node237_r & ~pixel[291];
      node246_r = node245_l & pixel[299];
      node246_l = node245_l & ~pixel[299];
      node247 = node246_l;
      node248 = node246_r;
      node249_r = node245_r & pixel[207];
      node249_l = node245_r & ~pixel[207];
      node250 = node249_l;
      node251 = node249_r;
      node252 = node220_r;
      node253_r = node219_r & pixel[355];
      node253_l = node219_r & ~pixel[355];
      node254_r = node253_l & pixel[382];
      node254_l = node253_l & ~pixel[382];
      node255_r = node254_l & pixel[235];
      node255_l = node254_l & ~pixel[235];
      node256_r = node255_l & pixel[380];
      node256_l = node255_l & ~pixel[380];
      node257_r = node256_l & pixel[570];
      node257_l = node256_l & ~pixel[570];
      node258 = node257_l;
      node259 = node257_r;
      node260_r = node256_r & pixel[573];
      node260_l = node256_r & ~pixel[573];
      node261 = node260_l;
      node262 = node260_r;
      node263_r = node255_r & pixel[681];
      node263_l = node255_r & ~pixel[681];
      node264_r = node263_l & pixel[403];
      node264_l = node263_l & ~pixel[403];
      node265 = node264_l;
      node266 = node264_r;
      node267_r = node263_r & pixel[350];
      node267_l = node263_r & ~pixel[350];
      node268 = node267_l;
      node269 = node267_r;
      node270_r = node254_r & pixel[573];
      node270_l = node254_r & ~pixel[573];
      node271_r = node270_l & pixel[156];
      node271_l = node270_l & ~pixel[156];
      node272_r = node271_l & pixel[203];
      node272_l = node271_l & ~pixel[203];
      node273 = node272_l;
      node274 = node272_r;
      node275_r = node271_r & pixel[598];
      node275_l = node271_r & ~pixel[598];
      node276 = node275_l;
      node277 = node275_r;
      node278_r = node270_r & pixel[131];
      node278_l = node270_r & ~pixel[131];
      node279_r = node278_l & pixel[542];
      node279_l = node278_l & ~pixel[542];
      node280 = node279_l;
      node281 = node279_r;
      node282_r = node278_r & pixel[599];
      node282_l = node278_r & ~pixel[599];
      node283 = node282_l;
      node284 = node282_r;
      node285_r = node253_r & pixel[160];
      node285_l = node253_r & ~pixel[160];
      node286_r = node285_l & pixel[457];
      node286_l = node285_l & ~pixel[457];
      node287_r = node286_l & pixel[156];
      node287_l = node286_l & ~pixel[156];
      node288_r = node287_l & pixel[430];
      node288_l = node287_l & ~pixel[430];
      node289 = node288_l;
      node290 = node288_r;
      node291_r = node287_r & pixel[403];
      node291_l = node287_r & ~pixel[403];
      node292 = node291_l;
      node293 = node291_r;
      node294_r = node286_r & pixel[235];
      node294_l = node286_r & ~pixel[235];
      node295_r = node294_l & pixel[569];
      node295_l = node294_l & ~pixel[569];
      node296 = node295_l;
      node297 = node295_r;
      node298_r = node294_r & pixel[568];
      node298_l = node294_r & ~pixel[568];
      node299 = node298_l;
      node300 = node298_r;
      node301_r = node285_r & pixel[484];
      node301_l = node285_r & ~pixel[484];
      node302_r = node301_l & pixel[594];
      node302_l = node301_l & ~pixel[594];
      node303_r = node302_l & pixel[678];
      node303_l = node302_l & ~pixel[678];
      node304 = node303_l;
      node305 = node303_r;
      node306_r = node302_r & pixel[426];
      node306_l = node302_r & ~pixel[426];
      node307 = node306_l;
      node308 = node306_r;
      node309_r = node301_r & pixel[621];
      node309_l = node301_r & ~pixel[621];
      node310_r = node309_l & pixel[572];
      node310_l = node309_l & ~pixel[572];
      node311 = node310_l;
      node312 = node310_r;
      node313 = node309_r;
      node314_r = node218_r & pixel[567];
      node314_l = node218_r & ~pixel[567];
      node315_r = node314_l & pixel[236];
      node315_l = node314_l & ~pixel[236];
      node316_r = node315_l & pixel[72];
      node316_l = node315_l & ~pixel[72];
      node317_r = node316_l & pixel[324];
      node317_l = node316_l & ~pixel[324];
      node318_r = node317_l & pixel[242];
      node318_l = node317_l & ~pixel[242];
      node319_r = node318_l & pixel[131];
      node319_l = node318_l & ~pixel[131];
      node320 = node319_l;
      node321 = node319_r;
      node322_r = node318_r & pixel[327];
      node322_l = node318_r & ~pixel[327];
      node323 = node322_l;
      node324 = node322_r;
      node325_r = node317_r & pixel[633];
      node325_l = node317_r & ~pixel[633];
      node326 = node325_l;
      node327_r = node325_r & pixel[573];
      node327_l = node325_r & ~pixel[573];
      node328 = node327_l;
      node329 = node327_r;
      node330 = node316_r;
      node331_r = node315_r & pixel[298];
      node331_l = node315_r & ~pixel[298];
      node332_r = node331_l & pixel[257];
      node332_l = node331_l & ~pixel[257];
      node333_r = node332_l & pixel[594];
      node333_l = node332_l & ~pixel[594];
      node334_r = node333_l & pixel[244];
      node334_l = node333_l & ~pixel[244];
      node335 = node334_l;
      node336 = node334_r;
      node337 = node333_r;
      node338 = node332_r;
      node339_r = node331_r & pixel[440];
      node339_l = node331_r & ~pixel[440];
      node340_r = node339_l & pixel[380];
      node340_l = node339_l & ~pixel[380];
      node341_r = node340_l & pixel[238];
      node341_l = node340_l & ~pixel[238];
      node342 = node341_l;
      node343 = node341_r;
      node344 = node340_r;
      node345_r = node339_r & pixel[269];
      node345_l = node339_r & ~pixel[269];
      node346 = node345_l;
      node347 = node345_r;
      node348_r = node314_r & pixel[327];
      node348_l = node314_r & ~pixel[327];
      node349_r = node348_l & pixel[453];
      node349_l = node348_l & ~pixel[453];
      node350_r = node349_l & pixel[515];
      node350_l = node349_l & ~pixel[515];
      node351 = node350_l;
      node352 = node350_r;
      node353 = node349_r;
      node354_r = node348_r & pixel[294];
      node354_l = node348_r & ~pixel[294];
      node355 = node354_l;
      node356 = node354_r;
      node357_r = node1_r & pixel[517];
      node357_l = node1_r & ~pixel[517];
      node358_r = node357_l & pixel[491];
      node358_l = node357_l & ~pixel[491];
      node359_r = node358_l & pixel[460];
      node359_l = node358_l & ~pixel[460];
      node360_r = node359_l & pixel[398];
      node360_l = node359_l & ~pixel[398];
      node361_r = node360_l & pixel[401];
      node361_l = node360_l & ~pixel[401];
      node362_r = node361_l & pixel[324];
      node362_l = node361_l & ~pixel[324];
      node363_r = node362_l & pixel[414];
      node363_l = node362_l & ~pixel[414];
      node364_r = node363_l & pixel[429];
      node364_l = node363_l & ~pixel[429];
      node365 = node364_l;
      node366 = node364_r;
      node367_r = node363_r & pixel[659];
      node367_l = node363_r & ~pixel[659];
      node368 = node367_l;
      node369 = node367_r;
      node370_r = node362_r & pixel[290];
      node370_l = node362_r & ~pixel[290];
      node371_r = node370_l & pixel[213];
      node371_l = node370_l & ~pixel[213];
      node372 = node371_l;
      node373 = node371_r;
      node374_r = node370_r & pixel[241];
      node374_l = node370_r & ~pixel[241];
      node375 = node374_l;
      node376 = node374_r;
      node377_r = node361_r & pixel[214];
      node377_l = node361_r & ~pixel[214];
      node378_r = node377_l & pixel[376];
      node378_l = node377_l & ~pixel[376];
      node379_r = node378_l & pixel[148];
      node379_l = node378_l & ~pixel[148];
      node380 = node379_l;
      node381 = node379_r;
      node382_r = node378_r & pixel[519];
      node382_l = node378_r & ~pixel[519];
      node383 = node382_l;
      node384 = node382_r;
      node385_r = node377_r & pixel[434];
      node385_l = node377_r & ~pixel[434];
      node386_r = node385_l & pixel[688];
      node386_l = node385_l & ~pixel[688];
      node387 = node386_l;
      node388 = node386_r;
      node389_r = node385_r & pixel[513];
      node389_l = node385_r & ~pixel[513];
      node390 = node389_l;
      node391 = node389_r;
      node392_r = node360_r & pixel[722];
      node392_l = node360_r & ~pixel[722];
      node393_r = node392_l & pixel[330];
      node393_l = node392_l & ~pixel[330];
      node394_r = node393_l & pixel[511];
      node394_l = node393_l & ~pixel[511];
      node395_r = node394_l & pixel[453];
      node395_l = node394_l & ~pixel[453];
      node396 = node395_l;
      node397 = node395_r;
      node398_r = node394_r & pixel[426];
      node398_l = node394_r & ~pixel[426];
      node399 = node398_l;
      node400 = node398_r;
      node401_r = node393_r & pixel[102];
      node401_l = node393_r & ~pixel[102];
      node402_r = node401_l & pixel[629];
      node402_l = node401_l & ~pixel[629];
      node403 = node402_l;
      node404 = node402_r;
      node405_r = node401_r & pixel[407];
      node405_l = node401_r & ~pixel[407];
      node406 = node405_l;
      node407 = node405_r;
      node408 = node392_r;
      node409_r = node359_r & pixel[132];
      node409_l = node359_r & ~pixel[132];
      node410_r = node409_l & pixel[125];
      node410_l = node409_l & ~pixel[125];
      node411_r = node410_l & pixel[156];
      node411_l = node410_l & ~pixel[156];
      node412_r = node411_l & pixel[356];
      node412_l = node411_l & ~pixel[356];
      node413_r = node412_l & pixel[438];
      node413_l = node412_l & ~pixel[438];
      node414 = node413_l;
      node415 = node413_r;
      node416_r = node412_r & pixel[343];
      node416_l = node412_r & ~pixel[343];
      node417 = node416_l;
      node418 = node416_r;
      node419_r = node411_r & pixel[214];
      node419_l = node411_r & ~pixel[214];
      node420_r = node419_l & pixel[687];
      node420_l = node419_l & ~pixel[687];
      node421 = node420_l;
      node422 = node420_r;
      node423_r = node419_r & pixel[408];
      node423_l = node419_r & ~pixel[408];
      node424 = node423_l;
      node425 = node423_r;
      node426_r = node410_r & pixel[317];
      node426_l = node410_r & ~pixel[317];
      node427 = node426_l;
      node428_r = node426_r & pixel[436];
      node428_l = node426_r & ~pixel[436];
      node429_r = node428_l & pixel[147];
      node429_l = node428_l & ~pixel[147];
      node430 = node429_l;
      node431 = node429_r;
      node432_r = node428_r & pixel[182];
      node432_l = node428_r & ~pixel[182];
      node433 = node432_l;
      node434 = node432_r;
      node435_r = node409_r & pixel[654];
      node435_l = node409_r & ~pixel[654];
      node436_r = node435_l & pixel[663];
      node436_l = node435_l & ~pixel[663];
      node437_r = node436_l & pixel[600];
      node437_l = node436_l & ~pixel[600];
      node438_r = node437_l & pixel[105];
      node438_l = node437_l & ~pixel[105];
      node439 = node438_l;
      node440 = node438_r;
      node441_r = node437_r & pixel[455];
      node441_l = node437_r & ~pixel[455];
      node442 = node441_l;
      node443 = node441_r;
      node444_r = node436_r & pixel[515];
      node444_l = node436_r & ~pixel[515];
      node445 = node444_l;
      node446 = node444_r;
      node447_r = node435_r & pixel[206];
      node447_l = node435_r & ~pixel[206];
      node448_r = node447_l & pixel[409];
      node448_l = node447_l & ~pixel[409];
      node449_r = node448_l & pixel[623];
      node449_l = node448_l & ~pixel[623];
      node450 = node449_l;
      node451 = node449_r;
      node452_r = node448_r & pixel[514];
      node452_l = node448_r & ~pixel[514];
      node453 = node452_l;
      node454 = node452_r;
      node455 = node447_r;
      node456_r = node358_r & pixel[439];
      node456_l = node358_r & ~pixel[439];
      node457_r = node456_l & pixel[248];
      node457_l = node456_l & ~pixel[248];
      node458_r = node457_l & pixel[461];
      node458_l = node457_l & ~pixel[461];
      node459_r = node458_l & pixel[295];
      node459_l = node458_l & ~pixel[295];
      node460_r = node459_l & pixel[654];
      node460_l = node459_l & ~pixel[654];
      node461 = node460_l;
      node462_r = node460_r & pixel[270];
      node462_l = node460_r & ~pixel[270];
      node463 = node462_l;
      node464 = node462_r;
      node465_r = node459_r & pixel[96];
      node465_l = node459_r & ~pixel[96];
      node466_r = node465_l & pixel[402];
      node466_l = node465_l & ~pixel[402];
      node467 = node466_l;
      node468 = node466_r;
      node469 = node465_r;
      node470_r = node458_r & pixel[375];
      node470_l = node458_r & ~pixel[375];
      node471_r = node470_l & pixel[437];
      node471_l = node470_l & ~pixel[437];
      node472_r = node471_l & pixel[685];
      node472_l = node471_l & ~pixel[685];
      node473 = node472_l;
      node474 = node472_r;
      node475_r = node471_r & pixel[568];
      node475_l = node471_r & ~pixel[568];
      node476 = node475_l;
      node477 = node475_r;
      node478_r = node470_r & pixel[428];
      node478_l = node470_r & ~pixel[428];
      node479_r = node478_l & pixel[355];
      node479_l = node478_l & ~pixel[355];
      node480 = node479_l;
      node481 = node479_r;
      node482_r = node478_r & pixel[240];
      node482_l = node478_r & ~pixel[240];
      node483 = node482_l;
      node484 = node482_r;
      node485_r = node457_r & pixel[515];
      node485_l = node457_r & ~pixel[515];
      node486_r = node485_l & pixel[425];
      node486_l = node485_l & ~pixel[425];
      node487 = node486_l;
      node488 = node486_r;
      node489_r = node485_r & pixel[380];
      node489_l = node485_r & ~pixel[380];
      node490 = node489_l;
      node491 = node489_r;
      node492_r = node456_r & pixel[461];
      node492_l = node456_r & ~pixel[461];
      node493_r = node492_l & pixel[498];
      node493_l = node492_l & ~pixel[498];
      node494_r = node493_l & pixel[187];
      node494_l = node493_l & ~pixel[187];
      node495_r = node494_l & pixel[214];
      node495_l = node494_l & ~pixel[214];
      node496_r = node495_l & pixel[296];
      node496_l = node495_l & ~pixel[296];
      node497 = node496_l;
      node498 = node496_r;
      node499_r = node495_r & pixel[347];
      node499_l = node495_r & ~pixel[347];
      node500 = node499_l;
      node501 = node499_r;
      node502_r = node494_r & pixel[328];
      node502_l = node494_r & ~pixel[328];
      node503_r = node502_l & pixel[344];
      node503_l = node502_l & ~pixel[344];
      node504 = node503_l;
      node505 = node503_r;
      node506_r = node502_r & pixel[265];
      node506_l = node502_r & ~pixel[265];
      node507 = node506_l;
      node508 = node506_r;
      node509_r = node493_r & pixel[626];
      node509_l = node493_r & ~pixel[626];
      node510 = node509_l;
      node511_r = node509_r & pixel[657];
      node511_l = node509_r & ~pixel[657];
      node512_r = node511_l & pixel[317];
      node512_l = node511_l & ~pixel[317];
      node513 = node512_l;
      node514 = node512_r;
      node515 = node511_r;
      node516_r = node492_r & pixel[155];
      node516_l = node492_r & ~pixel[155];
      node517_r = node516_l & pixel[346];
      node517_l = node516_l & ~pixel[346];
      node518_r = node517_l & pixel[316];
      node518_l = node517_l & ~pixel[316];
      node519_r = node518_l & pixel[573];
      node519_l = node518_l & ~pixel[573];
      node520 = node519_l;
      node521 = node519_r;
      node522_r = node518_r & pixel[601];
      node522_l = node518_r & ~pixel[601];
      node523 = node522_l;
      node524 = node522_r;
      node525_r = node517_r & pixel[652];
      node525_l = node517_r & ~pixel[652];
      node526_r = node525_l & pixel[103];
      node526_l = node525_l & ~pixel[103];
      node527 = node526_l;
      node528 = node526_r;
      node529 = node525_r;
      node530_r = node516_r & pixel[373];
      node530_l = node516_r & ~pixel[373];
      node531_r = node530_l & pixel[484];
      node531_l = node530_l & ~pixel[484];
      node532_r = node531_l & pixel[678];
      node532_l = node531_l & ~pixel[678];
      node533 = node532_l;
      node534 = node532_r;
      node535_r = node531_r & pixel[237];
      node535_l = node531_r & ~pixel[237];
      node536 = node535_l;
      node537 = node535_r;
      node538_r = node530_r & pixel[597];
      node538_l = node530_r & ~pixel[597];
      node539_r = node538_l & pixel[372];
      node539_l = node538_l & ~pixel[372];
      node540 = node539_l;
      node541 = node539_r;
      node542_r = node538_r & pixel[272];
      node542_l = node538_r & ~pixel[272];
      node543 = node542_l;
      node544 = node542_r;
      node545_r = node357_r & pixel[359];
      node545_l = node357_r & ~pixel[359];
      node546_r = node545_l & pixel[347];
      node546_l = node545_l & ~pixel[347];
      node547_r = node546_l & pixel[343];
      node547_l = node546_l & ~pixel[343];
      node548_r = node547_l & pixel[249];
      node548_l = node547_l & ~pixel[249];
      node549_r = node548_l & pixel[687];
      node549_l = node548_l & ~pixel[687];
      node550_r = node549_l & pixel[317];
      node550_l = node549_l & ~pixel[317];
      node551_r = node550_l & pixel[154];
      node551_l = node550_l & ~pixel[154];
      node552 = node551_l;
      node553 = node551_r;
      node554_r = node550_r & pixel[440];
      node554_l = node550_r & ~pixel[440];
      node555 = node554_l;
      node556 = node554_r;
      node557_r = node549_r & pixel[229];
      node557_l = node549_r & ~pixel[229];
      node558_r = node557_l & pixel[548];
      node558_l = node557_l & ~pixel[548];
      node559 = node558_l;
      node560 = node558_r;
      node561 = node557_r;
      node562_r = node548_r & pixel[385];
      node562_l = node548_r & ~pixel[385];
      node563 = node562_l;
      node564 = node562_r;
      node565_r = node547_r & pixel[571];
      node565_l = node547_r & ~pixel[571];
      node566_r = node565_l & pixel[454];
      node566_l = node565_l & ~pixel[454];
      node567_r = node566_l & pixel[373];
      node567_l = node566_l & ~pixel[373];
      node568_r = node567_l & pixel[150];
      node568_l = node567_l & ~pixel[150];
      node569 = node568_l;
      node570 = node568_r;
      node571_r = node567_r & pixel[315];
      node571_l = node567_r & ~pixel[315];
      node572 = node571_l;
      node573 = node571_r;
      node574_r = node566_r & pixel[427];
      node574_l = node566_r & ~pixel[427];
      node575 = node574_l;
      node576_r = node574_r & pixel[267];
      node576_l = node574_r & ~pixel[267];
      node577 = node576_l;
      node578 = node576_r;
      node579_r = node565_r & pixel[242];
      node579_l = node565_r & ~pixel[242];
      node580_r = node579_l & pixel[470];
      node580_l = node579_l & ~pixel[470];
      node581_r = node580_l & pixel[297];
      node581_l = node580_l & ~pixel[297];
      node582 = node581_l;
      node583 = node581_r;
      node584_r = node580_r & pixel[431];
      node584_l = node580_r & ~pixel[431];
      node585 = node584_l;
      node586 = node584_r;
      node587_r = node579_r & pixel[441];
      node587_l = node579_r & ~pixel[441];
      node588_r = node587_l & pixel[135];
      node588_l = node587_l & ~pixel[135];
      node589 = node588_l;
      node590 = node588_r;
      node591_r = node587_r & pixel[666];
      node591_l = node587_r & ~pixel[666];
      node592 = node591_l;
      node593 = node591_r;
      node594_r = node546_r & pixel[300];
      node594_l = node546_r & ~pixel[300];
      node595_r = node594_l & pixel[456];
      node595_l = node594_l & ~pixel[456];
      node596_r = node595_l & pixel[408];
      node596_l = node595_l & ~pixel[408];
      node597_r = node596_l & pixel[131];
      node597_l = node596_l & ~pixel[131];
      node598_r = node597_l & pixel[97];
      node598_l = node597_l & ~pixel[97];
      node599 = node598_l;
      node600 = node598_r;
      node601_r = node597_r & pixel[262];
      node601_l = node597_r & ~pixel[262];
      node602 = node601_l;
      node603 = node601_r;
      node604_r = node596_r & pixel[520];
      node604_l = node596_r & ~pixel[520];
      node605_r = node604_l & pixel[549];
      node605_l = node604_l & ~pixel[549];
      node606 = node605_l;
      node607 = node605_r;
      node608_r = node604_r & pixel[622];
      node608_l = node604_r & ~pixel[622];
      node609 = node608_l;
      node610 = node608_r;
      node611_r = node595_r & pixel[438];
      node611_l = node595_r & ~pixel[438];
      node612_r = node611_l & pixel[440];
      node612_l = node611_l & ~pixel[440];
      node613_r = node612_l & pixel[432];
      node613_l = node612_l & ~pixel[432];
      node614 = node613_l;
      node615 = node613_r;
      node616_r = node612_r & pixel[183];
      node616_l = node612_r & ~pixel[183];
      node617 = node616_l;
      node618 = node616_r;
      node619_r = node611_r & pixel[550];
      node619_l = node611_r & ~pixel[550];
      node620_r = node619_l & pixel[569];
      node620_l = node619_l & ~pixel[569];
      node621 = node620_l;
      node622 = node620_r;
      node623_r = node619_r & pixel[440];
      node623_l = node619_r & ~pixel[440];
      node624 = node623_l;
      node625 = node623_r;
      node626_r = node594_r & pixel[465];
      node626_l = node594_r & ~pixel[465];
      node627_r = node626_l & pixel[382];
      node627_l = node626_l & ~pixel[382];
      node628_r = node627_l & pixel[496];
      node628_l = node627_l & ~pixel[496];
      node629_r = node628_l & pixel[100];
      node629_l = node628_l & ~pixel[100];
      node630 = node629_l;
      node631 = node629_r;
      node632_r = node628_r & pixel[468];
      node632_l = node628_r & ~pixel[468];
      node633 = node632_l;
      node634 = node632_r;
      node635_r = node627_r & pixel[405];
      node635_l = node627_r & ~pixel[405];
      node636_r = node635_l & pixel[495];
      node636_l = node635_l & ~pixel[495];
      node637 = node636_l;
      node638 = node636_r;
      node639_r = node635_r & pixel[653];
      node639_l = node635_r & ~pixel[653];
      node640 = node639_l;
      node641 = node639_r;
      node642_r = node626_r & pixel[407];
      node642_l = node626_r & ~pixel[407];
      node643_r = node642_l & pixel[488];
      node643_l = node642_l & ~pixel[488];
      node644_r = node643_l & pixel[600];
      node644_l = node643_l & ~pixel[600];
      node645 = node644_l;
      node646 = node644_r;
      node647_r = node643_r & pixel[569];
      node647_l = node643_r & ~pixel[569];
      node648 = node647_l;
      node649 = node647_r;
      node650_r = node642_r & pixel[426];
      node650_l = node642_r & ~pixel[426];
      node651_r = node650_l & pixel[403];
      node651_l = node650_l & ~pixel[403];
      node652 = node651_l;
      node653 = node651_r;
      node654_r = node650_r & pixel[131];
      node654_l = node650_r & ~pixel[131];
      node655 = node654_l;
      node656 = node654_r;
      node657_r = node545_r & pixel[426];
      node657_l = node545_r & ~pixel[426];
      node658_r = node657_l & pixel[408];
      node658_l = node657_l & ~pixel[408];
      node659_r = node658_l & pixel[376];
      node659_l = node658_l & ~pixel[376];
      node660_r = node659_l & pixel[439];
      node660_l = node659_l & ~pixel[439];
      node661_r = node660_l & pixel[607];
      node661_l = node660_l & ~pixel[607];
      node662 = node661_l;
      node663 = node661_r;
      node664_r = node660_r & pixel[344];
      node664_l = node660_r & ~pixel[344];
      node665_r = node664_l & pixel[320];
      node665_l = node664_l & ~pixel[320];
      node666 = node665_l;
      node667 = node665_r;
      node668 = node664_r;
      node669_r = node659_r & pixel[626];
      node669_l = node659_r & ~pixel[626];
      node670_r = node669_l & pixel[440];
      node670_l = node669_l & ~pixel[440];
      node671 = node670_l;
      node672 = node670_r;
      node673_r = node669_r & pixel[442];
      node673_l = node669_r & ~pixel[442];
      node674_r = node673_l & pixel[384];
      node674_l = node673_l & ~pixel[384];
      node675 = node674_l;
      node676 = node674_r;
      node677 = node673_r;
      node678_r = node658_r & pixel[521];
      node678_l = node658_r & ~pixel[521];
      node679_r = node678_l & pixel[523];
      node679_l = node678_l & ~pixel[523];
      node680_r = node679_l & pixel[494];
      node680_l = node679_l & ~pixel[494];
      node681_r = node680_l & pixel[431];
      node681_l = node680_l & ~pixel[431];
      node682 = node681_l;
      node683 = node681_r;
      node684_r = node680_r & pixel[375];
      node684_l = node680_r & ~pixel[375];
      node685 = node684_l;
      node686 = node684_r;
      node687_r = node679_r & pixel[660];
      node687_l = node679_r & ~pixel[660];
      node688 = node687_l;
      node689 = node687_r;
      node690_r = node678_r & pixel[374];
      node690_l = node678_r & ~pixel[374];
      node691 = node690_l;
      node692_r = node690_r & pixel[269];
      node692_l = node690_r & ~pixel[269];
      node693 = node692_l;
      node694 = node692_r;
      node695_r = node657_r & pixel[267];
      node695_l = node657_r & ~pixel[267];
      node696_r = node695_l & pixel[187];
      node696_l = node695_l & ~pixel[187];
      node697_r = node696_l & pixel[410];
      node697_l = node696_l & ~pixel[410];
      node698_r = node697_l & pixel[353];
      node698_l = node697_l & ~pixel[353];
      node699_r = node698_l & pixel[127];
      node699_l = node698_l & ~pixel[127];
      node700 = node699_l;
      node701 = node699_r;
      node702 = node698_r;
      node703_r = node697_r & pixel[270];
      node703_l = node697_r & ~pixel[270];
      node704_r = node703_l & pixel[634];
      node704_l = node703_l & ~pixel[634];
      node705 = node704_l;
      node706 = node704_r;
      node707_r = node703_r & pixel[431];
      node707_l = node703_r & ~pixel[431];
      node708 = node707_l;
      node709 = node707_r;
      node710_r = node696_r & pixel[461];
      node710_l = node696_r & ~pixel[461];
      node711 = node710_l;
      node712_r = node710_r & pixel[464];
      node712_l = node710_r & ~pixel[464];
      node713 = node712_l;
      node714_r = node712_r & pixel[232];
      node714_l = node712_r & ~pixel[232];
      node715 = node714_l;
      node716 = node714_r;
      node717_r = node695_r & pixel[690];
      node717_l = node695_r & ~pixel[690];
      node718_r = node717_l & pixel[77];
      node718_l = node717_l & ~pixel[77];
      node719_r = node718_l & pixel[435];
      node719_l = node718_l & ~pixel[435];
      node720_r = node719_l & pixel[265];
      node720_l = node719_l & ~pixel[265];
      node721 = node720_l;
      node722 = node720_r;
      node723_r = node719_r & pixel[299];
      node723_l = node719_r & ~pixel[299];
      node724 = node723_l;
      node725 = node723_r;
      node726 = node718_r;
      node727_r = node717_r & pixel[402];
      node727_l = node717_r & ~pixel[402];
      node728 = node727_l;
      node729 = node727_r;
      node730_r = node0_r & pixel[291];
      node730_l = node0_r & ~pixel[291];
      node731_r = node730_l & pixel[550];
      node731_l = node730_l & ~pixel[550];
      node732_r = node731_l & pixel[207];
      node732_l = node731_l & ~pixel[207];
      node733_r = node732_l & pixel[439];
      node733_l = node732_l & ~pixel[439];
      node734_r = node733_l & pixel[489];
      node734_l = node733_l & ~pixel[489];
      node735_r = node734_l & pixel[653];
      node735_l = node734_l & ~pixel[653];
      node736_r = node735_l & pixel[275];
      node736_l = node735_l & ~pixel[275];
      node737_r = node736_l & pixel[344];
      node737_l = node736_l & ~pixel[344];
      node738_r = node737_l & pixel[570];
      node738_l = node737_l & ~pixel[570];
      node739 = node738_l;
      node740 = node738_r;
      node741_r = node737_r & pixel[609];
      node741_l = node737_r & ~pixel[609];
      node742 = node741_l;
      node743 = node741_r;
      node744_r = node736_r & pixel[343];
      node744_l = node736_r & ~pixel[343];
      node745_r = node744_l & pixel[443];
      node745_l = node744_l & ~pixel[443];
      node746 = node745_l;
      node747 = node745_r;
      node748_r = node744_r & pixel[429];
      node748_l = node744_r & ~pixel[429];
      node749 = node748_l;
      node750 = node748_r;
      node751_r = node735_r & pixel[540];
      node751_l = node735_r & ~pixel[540];
      node752_r = node751_l & pixel[155];
      node752_l = node751_l & ~pixel[155];
      node753_r = node752_l & pixel[492];
      node753_l = node752_l & ~pixel[492];
      node754 = node753_l;
      node755 = node753_r;
      node756_r = node752_r & pixel[456];
      node756_l = node752_r & ~pixel[456];
      node757 = node756_l;
      node758 = node756_r;
      node759_r = node751_r & pixel[122];
      node759_l = node751_r & ~pixel[122];
      node760_r = node759_l & pixel[300];
      node760_l = node759_l & ~pixel[300];
      node761 = node760_l;
      node762 = node760_r;
      node763_r = node759_r & pixel[156];
      node763_l = node759_r & ~pixel[156];
      node764 = node763_l;
      node765 = node763_r;
      node766_r = node734_r & pixel[299];
      node766_l = node734_r & ~pixel[299];
      node767_r = node766_l & pixel[123];
      node767_l = node766_l & ~pixel[123];
      node768_r = node767_l & pixel[329];
      node768_l = node767_l & ~pixel[329];
      node769_r = node768_l & pixel[538];
      node769_l = node768_l & ~pixel[538];
      node770 = node769_l;
      node771 = node769_r;
      node772_r = node768_r & pixel[410];
      node772_l = node768_r & ~pixel[410];
      node773 = node772_l;
      node774 = node772_r;
      node775_r = node767_r & pixel[208];
      node775_l = node767_r & ~pixel[208];
      node776_r = node775_l & pixel[343];
      node776_l = node775_l & ~pixel[343];
      node777 = node776_l;
      node778 = node776_r;
      node779_r = node775_r & pixel[184];
      node779_l = node775_r & ~pixel[184];
      node780 = node779_l;
      node781 = node779_r;
      node782_r = node766_r & pixel[155];
      node782_l = node766_r & ~pixel[155];
      node783_r = node782_l & pixel[296];
      node783_l = node782_l & ~pixel[296];
      node784_r = node783_l & pixel[186];
      node784_l = node783_l & ~pixel[186];
      node785 = node784_l;
      node786 = node784_r;
      node787_r = node783_r & pixel[511];
      node787_l = node783_r & ~pixel[511];
      node788 = node787_l;
      node789 = node787_r;
      node790_r = node782_r & pixel[100];
      node790_l = node782_r & ~pixel[100];
      node791_r = node790_l & pixel[513];
      node791_l = node790_l & ~pixel[513];
      node792 = node791_l;
      node793 = node791_r;
      node794_r = node790_r & pixel[598];
      node794_l = node790_r & ~pixel[598];
      node795 = node794_l;
      node796 = node794_r;
      node797_r = node733_r & pixel[567];
      node797_l = node733_r & ~pixel[567];
      node798_r = node797_l & pixel[454];
      node798_l = node797_l & ~pixel[454];
      node799_r = node798_l & pixel[488];
      node799_l = node798_l & ~pixel[488];
      node800_r = node799_l & pixel[463];
      node800_l = node799_l & ~pixel[463];
      node801_r = node800_l & pixel[486];
      node801_l = node800_l & ~pixel[486];
      node802 = node801_l;
      node803 = node801_r;
      node804_r = node800_r & pixel[541];
      node804_l = node800_r & ~pixel[541];
      node805 = node804_l;
      node806 = node804_r;
      node807_r = node799_r & pixel[549];
      node807_l = node799_r & ~pixel[549];
      node808_r = node807_l & pixel[429];
      node808_l = node807_l & ~pixel[429];
      node809 = node808_l;
      node810 = node808_r;
      node811_r = node807_r & pixel[231];
      node811_l = node807_r & ~pixel[231];
      node812 = node811_l;
      node813 = node811_r;
      node814_r = node798_r & pixel[316];
      node814_l = node798_r & ~pixel[316];
      node815_r = node814_l & pixel[657];
      node815_l = node814_l & ~pixel[657];
      node816_r = node815_l & pixel[263];
      node816_l = node815_l & ~pixel[263];
      node817 = node816_l;
      node818 = node816_r;
      node819_r = node815_r & pixel[209];
      node819_l = node815_r & ~pixel[209];
      node820 = node819_l;
      node821 = node819_r;
      node822 = node814_r;
      node823_r = node797_r & pixel[488];
      node823_l = node797_r & ~pixel[488];
      node824_r = node823_l & pixel[294];
      node824_l = node823_l & ~pixel[294];
      node825_r = node824_l & pixel[381];
      node825_l = node824_l & ~pixel[381];
      node826 = node825_l;
      node827_r = node825_r & pixel[464];
      node827_l = node825_r & ~pixel[464];
      node828 = node827_l;
      node829 = node827_r;
      node830_r = node824_r & pixel[430];
      node830_l = node824_r & ~pixel[430];
      node831_r = node830_l & pixel[543];
      node831_l = node830_l & ~pixel[543];
      node832 = node831_l;
      node833 = node831_r;
      node834_r = node830_r & pixel[636];
      node834_l = node830_r & ~pixel[636];
      node835 = node834_l;
      node836 = node834_r;
      node837_r = node823_r & pixel[469];
      node837_l = node823_r & ~pixel[469];
      node838_r = node837_l & pixel[407];
      node838_l = node837_l & ~pixel[407];
      node839 = node838_l;
      node840_r = node838_r & pixel[521];
      node840_l = node838_r & ~pixel[521];
      node841 = node840_l;
      node842 = node840_r;
      node843_r = node837_r & pixel[320];
      node843_l = node837_r & ~pixel[320];
      node844_r = node843_l & pixel[318];
      node844_l = node843_l & ~pixel[318];
      node845 = node844_l;
      node846 = node844_r;
      node847_r = node843_r & pixel[436];
      node847_l = node843_r & ~pixel[436];
      node848 = node847_l;
      node849 = node847_r;
      node850_r = node732_r & pixel[515];
      node850_l = node732_r & ~pixel[515];
      node851_r = node850_l & pixel[553];
      node851_l = node850_l & ~pixel[553];
      node852_r = node851_l & pixel[317];
      node852_l = node851_l & ~pixel[317];
      node853_r = node852_l & pixel[652];
      node853_l = node852_l & ~pixel[652];
      node854_r = node853_l & pixel[261];
      node854_l = node853_l & ~pixel[261];
      node855_r = node854_l & pixel[321];
      node855_l = node854_l & ~pixel[321];
      node856 = node855_l;
      node857 = node855_r;
      node858_r = node854_r & pixel[491];
      node858_l = node854_r & ~pixel[491];
      node859 = node858_l;
      node860 = node858_r;
      node861_r = node853_r & pixel[412];
      node861_l = node853_r & ~pixel[412];
      node862_r = node861_l & pixel[454];
      node862_l = node861_l & ~pixel[454];
      node863 = node862_l;
      node864 = node862_r;
      node865_r = node861_r & pixel[598];
      node865_l = node861_r & ~pixel[598];
      node866 = node865_l;
      node867 = node865_r;
      node868_r = node852_r & pixel[208];
      node868_l = node852_r & ~pixel[208];
      node869_r = node868_l & pixel[154];
      node869_l = node868_l & ~pixel[154];
      node870 = node869_l;
      node871_r = node869_r & pixel[600];
      node871_l = node869_r & ~pixel[600];
      node872 = node871_l;
      node873 = node871_r;
      node874_r = node868_r & pixel[156];
      node874_l = node868_r & ~pixel[156];
      node875_r = node874_l & pixel[159];
      node875_l = node874_l & ~pixel[159];
      node876 = node875_l;
      node877 = node875_r;
      node878_r = node874_r & pixel[407];
      node878_l = node874_r & ~pixel[407];
      node879 = node878_l;
      node880 = node878_r;
      node881_r = node851_r & pixel[174];
      node881_l = node851_r & ~pixel[174];
      node882_r = node881_l & pixel[288];
      node882_l = node881_l & ~pixel[288];
      node883_r = node882_l & pixel[342];
      node883_l = node882_l & ~pixel[342];
      node884_r = node883_l & pixel[546];
      node884_l = node883_l & ~pixel[546];
      node885 = node884_l;
      node886 = node884_r;
      node887_r = node883_r & pixel[297];
      node887_l = node883_r & ~pixel[297];
      node888 = node887_l;
      node889 = node887_r;
      node890_r = node882_r & pixel[270];
      node890_l = node882_r & ~pixel[270];
      node891_r = node890_l & pixel[271];
      node891_l = node890_l & ~pixel[271];
      node892 = node891_l;
      node893 = node891_r;
      node894_r = node890_r & pixel[297];
      node894_l = node890_r & ~pixel[297];
      node895 = node894_l;
      node896 = node894_r;
      node897_r = node881_r & pixel[345];
      node897_l = node881_r & ~pixel[345];
      node898_r = node897_l & pixel[173];
      node898_l = node897_l & ~pixel[173];
      node899_r = node898_l & pixel[205];
      node899_l = node898_l & ~pixel[205];
      node900 = node899_l;
      node901 = node899_r;
      node902 = node898_r;
      node903_r = node897_r & pixel[186];
      node903_l = node897_r & ~pixel[186];
      node904_r = node903_l & pixel[267];
      node904_l = node903_l & ~pixel[267];
      node905 = node904_l;
      node906 = node904_r;
      node907_r = node903_r & pixel[296];
      node907_l = node903_r & ~pixel[296];
      node908 = node907_l;
      node909 = node907_r;
      node910_r = node850_r & pixel[127];
      node910_l = node850_r & ~pixel[127];
      node911_r = node910_l & pixel[150];
      node911_l = node910_l & ~pixel[150];
      node912_r = node911_l & pixel[432];
      node912_l = node911_l & ~pixel[432];
      node913_r = node912_l & pixel[320];
      node913_l = node912_l & ~pixel[320];
      node914_r = node913_l & pixel[240];
      node914_l = node913_l & ~pixel[240];
      node915 = node914_l;
      node916 = node914_r;
      node917_r = node913_r & pixel[155];
      node917_l = node913_r & ~pixel[155];
      node918 = node917_l;
      node919 = node917_r;
      node920_r = node912_r & pixel[627];
      node920_l = node912_r & ~pixel[627];
      node921_r = node920_l & pixel[345];
      node921_l = node920_l & ~pixel[345];
      node922 = node921_l;
      node923 = node921_r;
      node924_r = node920_r & pixel[157];
      node924_l = node920_r & ~pixel[157];
      node925 = node924_l;
      node926 = node924_r;
      node927_r = node911_r & pixel[374];
      node927_l = node911_r & ~pixel[374];
      node928_r = node927_l & pixel[679];
      node928_l = node927_l & ~pixel[679];
      node929_r = node928_l & pixel[682];
      node929_l = node928_l & ~pixel[682];
      node930 = node929_l;
      node931 = node929_r;
      node932_r = node928_r & pixel[258];
      node932_l = node928_r & ~pixel[258];
      node933 = node932_l;
      node934 = node932_r;
      node935_r = node927_r & pixel[285];
      node935_l = node927_r & ~pixel[285];
      node936_r = node935_l & pixel[581];
      node936_l = node935_l & ~pixel[581];
      node937 = node936_l;
      node938 = node936_r;
      node939 = node935_r;
      node940_r = node910_r & pixel[314];
      node940_l = node910_r & ~pixel[314];
      node941_r = node940_l & pixel[356];
      node941_l = node940_l & ~pixel[356];
      node942_r = node941_l & pixel[270];
      node942_l = node941_l & ~pixel[270];
      node943_r = node942_l & pixel[659];
      node943_l = node942_l & ~pixel[659];
      node944 = node943_l;
      node945 = node943_r;
      node946_r = node942_r & pixel[346];
      node946_l = node942_r & ~pixel[346];
      node947 = node946_l;
      node948 = node946_r;
      node949_r = node941_r & pixel[151];
      node949_l = node941_r & ~pixel[151];
      node950 = node949_l;
      node951_r = node949_r & pixel[330];
      node951_l = node949_r & ~pixel[330];
      node952 = node951_l;
      node953 = node951_r;
      node954_r = node940_r & pixel[539];
      node954_l = node940_r & ~pixel[539];
      node955_r = node954_l & pixel[181];
      node955_l = node954_l & ~pixel[181];
      node956 = node955_l;
      node957_r = node955_r & pixel[217];
      node957_l = node955_r & ~pixel[217];
      node958 = node957_l;
      node959 = node957_r;
      node960 = node954_r;
      node961_r = node731_r & pixel[653];
      node961_l = node731_r & ~pixel[653];
      node962_r = node961_l & pixel[438];
      node962_l = node961_l & ~pixel[438];
      node963_r = node962_l & pixel[386];
      node963_l = node962_l & ~pixel[386];
      node964_r = node963_l & pixel[345];
      node964_l = node963_l & ~pixel[345];
      node965_r = node964_l & pixel[572];
      node965_l = node964_l & ~pixel[572];
      node966_r = node965_l & pixel[657];
      node966_l = node965_l & ~pixel[657];
      node967_r = node966_l & pixel[542];
      node967_l = node966_l & ~pixel[542];
      node968 = node967_l;
      node969 = node967_r;
      node970_r = node966_r & pixel[515];
      node970_l = node966_r & ~pixel[515];
      node971 = node970_l;
      node972 = node970_r;
      node973_r = node965_r & pixel[540];
      node973_l = node965_r & ~pixel[540];
      node974_r = node973_l & pixel[217];
      node974_l = node973_l & ~pixel[217];
      node975 = node974_l;
      node976 = node974_r;
      node977_r = node973_r & pixel[554];
      node977_l = node973_r & ~pixel[554];
      node978 = node977_l;
      node979 = node977_r;
      node980_r = node964_r & pixel[633];
      node980_l = node964_r & ~pixel[633];
      node981_r = node980_l & pixel[267];
      node981_l = node980_l & ~pixel[267];
      node982_r = node981_l & pixel[289];
      node982_l = node981_l & ~pixel[289];
      node983 = node982_l;
      node984 = node982_r;
      node985_r = node981_r & pixel[230];
      node985_l = node981_r & ~pixel[230];
      node986 = node985_l;
      node987 = node985_r;
      node988_r = node980_r & pixel[299];
      node988_l = node980_r & ~pixel[299];
      node989_r = node988_l & pixel[573];
      node989_l = node988_l & ~pixel[573];
      node990 = node989_l;
      node991 = node989_r;
      node992_r = node988_r & pixel[316];
      node992_l = node988_r & ~pixel[316];
      node993 = node992_l;
      node994 = node992_r;
      node995_r = node963_r & pixel[182];
      node995_l = node963_r & ~pixel[182];
      node996_r = node995_l & pixel[103];
      node996_l = node995_l & ~pixel[103];
      node997_r = node996_l & pixel[238];
      node997_l = node996_l & ~pixel[238];
      node998_r = node997_l & pixel[320];
      node998_l = node997_l & ~pixel[320];
      node999 = node998_l;
      node1000 = node998_r;
      node1001_r = node997_r & pixel[382];
      node1001_l = node997_r & ~pixel[382];
      node1002 = node1001_l;
      node1003 = node1001_r;
      node1004_r = node996_r & pixel[428];
      node1004_l = node996_r & ~pixel[428];
      node1005 = node1004_l;
      node1006 = node1004_r;
      node1007_r = node995_r & pixel[316];
      node1007_l = node995_r & ~pixel[316];
      node1008_r = node1007_l & pixel[602];
      node1008_l = node1007_l & ~pixel[602];
      node1009 = node1008_l;
      node1010_r = node1008_r & pixel[325];
      node1010_l = node1008_r & ~pixel[325];
      node1011 = node1010_l;
      node1012 = node1010_r;
      node1013_r = node1007_r & pixel[685];
      node1013_l = node1007_r & ~pixel[685];
      node1014_r = node1013_l & pixel[548];
      node1014_l = node1013_l & ~pixel[548];
      node1015 = node1014_l;
      node1016 = node1014_r;
      node1017_r = node1013_r & pixel[541];
      node1017_l = node1013_r & ~pixel[541];
      node1018 = node1017_l;
      node1019 = node1017_r;
      node1020_r = node962_r & pixel[597];
      node1020_l = node962_r & ~pixel[597];
      node1021_r = node1020_l & pixel[211];
      node1021_l = node1020_l & ~pixel[211];
      node1022_r = node1021_l & pixel[498];
      node1022_l = node1021_l & ~pixel[498];
      node1023_r = node1022_l & pixel[293];
      node1023_l = node1022_l & ~pixel[293];
      node1024_r = node1023_l & pixel[427];
      node1024_l = node1023_l & ~pixel[427];
      node1025 = node1024_l;
      node1026 = node1024_r;
      node1027_r = node1023_r & pixel[287];
      node1027_l = node1023_r & ~pixel[287];
      node1028 = node1027_l;
      node1029 = node1027_r;
      node1030_r = node1022_r & pixel[662];
      node1030_l = node1022_r & ~pixel[662];
      node1031_r = node1030_l & pixel[542];
      node1031_l = node1030_l & ~pixel[542];
      node1032 = node1031_l;
      node1033 = node1031_r;
      node1034_r = node1030_r & pixel[426];
      node1034_l = node1030_r & ~pixel[426];
      node1035 = node1034_l;
      node1036 = node1034_r;
      node1037_r = node1021_r & pixel[152];
      node1037_l = node1021_r & ~pixel[152];
      node1038_r = node1037_l & pixel[320];
      node1038_l = node1037_l & ~pixel[320];
      node1039_r = node1038_l & pixel[238];
      node1039_l = node1038_l & ~pixel[238];
      node1040 = node1039_l;
      node1041 = node1039_r;
      node1042_r = node1038_r & pixel[234];
      node1042_l = node1038_r & ~pixel[234];
      node1043 = node1042_l;
      node1044 = node1042_r;
      node1045_r = node1037_r & pixel[343];
      node1045_l = node1037_r & ~pixel[343];
      node1046_r = node1045_l & pixel[289];
      node1046_l = node1045_l & ~pixel[289];
      node1047 = node1046_l;
      node1048 = node1046_r;
      node1049_r = node1045_r & pixel[601];
      node1049_l = node1045_r & ~pixel[601];
      node1050 = node1049_l;
      node1051 = node1049_r;
      node1052_r = node1020_r & pixel[432];
      node1052_l = node1020_r & ~pixel[432];
      node1053_r = node1052_l & pixel[315];
      node1053_l = node1052_l & ~pixel[315];
      node1054_r = node1053_l & pixel[352];
      node1054_l = node1053_l & ~pixel[352];
      node1055_r = node1054_l & pixel[370];
      node1055_l = node1054_l & ~pixel[370];
      node1056 = node1055_l;
      node1057 = node1055_r;
      node1058_r = node1054_r & pixel[316];
      node1058_l = node1054_r & ~pixel[316];
      node1059 = node1058_l;
      node1060 = node1058_r;
      node1061_r = node1053_r & pixel[327];
      node1061_l = node1053_r & ~pixel[327];
      node1062_r = node1061_l & pixel[489];
      node1062_l = node1061_l & ~pixel[489];
      node1063 = node1062_l;
      node1064 = node1062_r;
      node1065_r = node1061_r & pixel[398];
      node1065_l = node1061_r & ~pixel[398];
      node1066 = node1065_l;
      node1067 = node1065_r;
      node1068_r = node1052_r & pixel[181];
      node1068_l = node1052_r & ~pixel[181];
      node1069_r = node1068_l & pixel[126];
      node1069_l = node1068_l & ~pixel[126];
      node1070_r = node1069_l & pixel[263];
      node1070_l = node1069_l & ~pixel[263];
      node1071 = node1070_l;
      node1072 = node1070_r;
      node1073_r = node1069_r & pixel[577];
      node1073_l = node1069_r & ~pixel[577];
      node1074 = node1073_l;
      node1075 = node1073_r;
      node1076_r = node1068_r & pixel[631];
      node1076_l = node1068_r & ~pixel[631];
      node1077_r = node1076_l & pixel[484];
      node1077_l = node1076_l & ~pixel[484];
      node1078 = node1077_l;
      node1079 = node1077_r;
      node1080_r = node1076_r & pixel[344];
      node1080_l = node1076_r & ~pixel[344];
      node1081 = node1080_l;
      node1082 = node1080_r;
      node1083_r = node961_r & pixel[541];
      node1083_l = node961_r & ~pixel[541];
      node1084_r = node1083_l & pixel[324];
      node1084_l = node1083_l & ~pixel[324];
      node1085_r = node1084_l & pixel[289];
      node1085_l = node1084_l & ~pixel[289];
      node1086_r = node1085_l & pixel[632];
      node1086_l = node1085_l & ~pixel[632];
      node1087_r = node1086_l & pixel[400];
      node1087_l = node1086_l & ~pixel[400];
      node1088_r = node1087_l & pixel[190];
      node1088_l = node1087_l & ~pixel[190];
      node1089 = node1088_l;
      node1090 = node1088_r;
      node1091_r = node1087_r & pixel[510];
      node1091_l = node1087_r & ~pixel[510];
      node1092 = node1091_l;
      node1093 = node1091_r;
      node1094_r = node1086_r & pixel[267];
      node1094_l = node1086_r & ~pixel[267];
      node1095_r = node1094_l & pixel[355];
      node1095_l = node1094_l & ~pixel[355];
      node1096 = node1095_l;
      node1097 = node1095_r;
      node1098_r = node1094_r & pixel[542];
      node1098_l = node1094_r & ~pixel[542];
      node1099 = node1098_l;
      node1100 = node1098_r;
      node1101_r = node1085_r & pixel[347];
      node1101_l = node1085_r & ~pixel[347];
      node1102_r = node1101_l & pixel[650];
      node1102_l = node1101_l & ~pixel[650];
      node1103_r = node1102_l & pixel[271];
      node1103_l = node1102_l & ~pixel[271];
      node1104 = node1103_l;
      node1105 = node1103_r;
      node1106 = node1102_r;
      node1107_r = node1101_r & pixel[457];
      node1107_l = node1101_r & ~pixel[457];
      node1108_r = node1107_l & pixel[432];
      node1108_l = node1107_l & ~pixel[432];
      node1109 = node1108_l;
      node1110 = node1108_r;
      node1111_r = node1107_r & pixel[149];
      node1111_l = node1107_r & ~pixel[149];
      node1112 = node1111_l;
      node1113 = node1111_r;
      node1114_r = node1084_r & pixel[544];
      node1114_l = node1084_r & ~pixel[544];
      node1115_r = node1114_l & pixel[416];
      node1115_l = node1114_l & ~pixel[416];
      node1116_r = node1115_l & pixel[315];
      node1116_l = node1115_l & ~pixel[315];
      node1117_r = node1116_l & pixel[135];
      node1117_l = node1116_l & ~pixel[135];
      node1118 = node1117_l;
      node1119 = node1117_r;
      node1120_r = node1116_r & pixel[634];
      node1120_l = node1116_r & ~pixel[634];
      node1121 = node1120_l;
      node1122 = node1120_r;
      node1123_r = node1115_r & pixel[402];
      node1123_l = node1115_r & ~pixel[402];
      node1124 = node1123_l;
      node1125_r = node1123_r & pixel[635];
      node1125_l = node1123_r & ~pixel[635];
      node1126 = node1125_l;
      node1127 = node1125_r;
      node1128_r = node1114_r & pixel[375];
      node1128_l = node1114_r & ~pixel[375];
      node1129_r = node1128_l & pixel[465];
      node1129_l = node1128_l & ~pixel[465];
      node1130_r = node1129_l & pixel[470];
      node1130_l = node1129_l & ~pixel[470];
      node1131 = node1130_l;
      node1132 = node1130_r;
      node1133 = node1129_r;
      node1134_r = node1128_r & pixel[219];
      node1134_l = node1128_r & ~pixel[219];
      node1135_r = node1134_l & pixel[315];
      node1135_l = node1134_l & ~pixel[315];
      node1136 = node1135_l;
      node1137 = node1135_r;
      node1138 = node1134_r;
      node1139_r = node1083_r & pixel[573];
      node1139_l = node1083_r & ~pixel[573];
      node1140_r = node1139_l & pixel[288];
      node1140_l = node1139_l & ~pixel[288];
      node1141_r = node1140_l & pixel[151];
      node1141_l = node1140_l & ~pixel[151];
      node1142_r = node1141_l & pixel[377];
      node1142_l = node1141_l & ~pixel[377];
      node1143_r = node1142_l & pixel[152];
      node1143_l = node1142_l & ~pixel[152];
      node1144 = node1143_l;
      node1145 = node1143_r;
      node1146_r = node1142_r & pixel[152];
      node1146_l = node1142_r & ~pixel[152];
      node1147 = node1146_l;
      node1148 = node1146_r;
      node1149_r = node1141_r & pixel[461];
      node1149_l = node1141_r & ~pixel[461];
      node1150_r = node1149_l & pixel[317];
      node1150_l = node1149_l & ~pixel[317];
      node1151 = node1150_l;
      node1152 = node1150_r;
      node1153_r = node1149_r & pixel[574];
      node1153_l = node1149_r & ~pixel[574];
      node1154 = node1153_l;
      node1155 = node1153_r;
      node1156_r = node1140_r & pixel[514];
      node1156_l = node1140_r & ~pixel[514];
      node1157_r = node1156_l & pixel[238];
      node1157_l = node1156_l & ~pixel[238];
      node1158_r = node1157_l & pixel[570];
      node1158_l = node1157_l & ~pixel[570];
      node1159 = node1158_l;
      node1160 = node1158_r;
      node1161_r = node1157_r & pixel[511];
      node1161_l = node1157_r & ~pixel[511];
      node1162 = node1161_l;
      node1163 = node1161_r;
      node1164_r = node1156_r & pixel[206];
      node1164_l = node1156_r & ~pixel[206];
      node1165_r = node1164_l & pixel[294];
      node1165_l = node1164_l & ~pixel[294];
      node1166 = node1165_l;
      node1167 = node1165_r;
      node1168_r = node1164_r & pixel[406];
      node1168_l = node1164_r & ~pixel[406];
      node1169 = node1168_l;
      node1170 = node1168_r;
      node1171_r = node1139_r & pixel[461];
      node1171_l = node1139_r & ~pixel[461];
      node1172_r = node1171_l & pixel[352];
      node1172_l = node1171_l & ~pixel[352];
      node1173_r = node1172_l & pixel[580];
      node1173_l = node1172_l & ~pixel[580];
      node1174_r = node1173_l & pixel[243];
      node1174_l = node1173_l & ~pixel[243];
      node1175 = node1174_l;
      node1176 = node1174_r;
      node1177 = node1173_r;
      node1178_r = node1172_r & pixel[487];
      node1178_l = node1172_r & ~pixel[487];
      node1179_r = node1178_l & pixel[270];
      node1179_l = node1178_l & ~pixel[270];
      node1180 = node1179_l;
      node1181 = node1179_r;
      node1182_r = node1178_r & pixel[383];
      node1182_l = node1178_r & ~pixel[383];
      node1183 = node1182_l;
      node1184 = node1182_r;
      node1185_r = node1171_r & pixel[438];
      node1185_l = node1171_r & ~pixel[438];
      node1186_r = node1185_l & pixel[266];
      node1186_l = node1185_l & ~pixel[266];
      node1187_r = node1186_l & pixel[357];
      node1187_l = node1186_l & ~pixel[357];
      node1188 = node1187_l;
      node1189 = node1187_r;
      node1190_r = node1186_r & pixel[487];
      node1190_l = node1186_r & ~pixel[487];
      node1191 = node1190_l;
      node1192 = node1190_r;
      node1193_r = node1185_r & pixel[323];
      node1193_l = node1185_r & ~pixel[323];
      node1194_r = node1193_l & pixel[552];
      node1194_l = node1193_l & ~pixel[552];
      node1195 = node1194_l;
      node1196 = node1194_r;
      node1197_r = node1193_r & pixel[486];
      node1197_l = node1193_r & ~pixel[486];
      node1198 = node1197_l;
      node1199 = node1197_r;
      node1200_r = node730_r & pixel[570];
      node1200_l = node730_r & ~pixel[570];
      node1201_r = node1200_l & pixel[597];
      node1201_l = node1200_l & ~pixel[597];
      node1202_r = node1201_l & pixel[297];
      node1202_l = node1201_l & ~pixel[297];
      node1203_r = node1202_l & pixel[515];
      node1203_l = node1202_l & ~pixel[515];
      node1204_r = node1203_l & pixel[546];
      node1204_l = node1203_l & ~pixel[546];
      node1205_r = node1204_l & pixel[184];
      node1205_l = node1204_l & ~pixel[184];
      node1206_r = node1205_l & pixel[327];
      node1206_l = node1205_l & ~pixel[327];
      node1207_r = node1206_l & pixel[520];
      node1207_l = node1206_l & ~pixel[520];
      node1208 = node1207_l;
      node1209 = node1207_r;
      node1210_r = node1206_r & pixel[239];
      node1210_l = node1206_r & ~pixel[239];
      node1211 = node1210_l;
      node1212 = node1210_r;
      node1213_r = node1205_r & pixel[345];
      node1213_l = node1205_r & ~pixel[345];
      node1214_r = node1213_l & pixel[329];
      node1214_l = node1213_l & ~pixel[329];
      node1215 = node1214_l;
      node1216 = node1214_r;
      node1217_r = node1213_r & pixel[294];
      node1217_l = node1213_r & ~pixel[294];
      node1218 = node1217_l;
      node1219 = node1217_r;
      node1220_r = node1204_r & pixel[212];
      node1220_l = node1204_r & ~pixel[212];
      node1221_r = node1220_l & pixel[353];
      node1221_l = node1220_l & ~pixel[353];
      node1222_r = node1221_l & pixel[382];
      node1222_l = node1221_l & ~pixel[382];
      node1223 = node1222_l;
      node1224 = node1222_r;
      node1225_r = node1221_r & pixel[268];
      node1225_l = node1221_r & ~pixel[268];
      node1226 = node1225_l;
      node1227 = node1225_r;
      node1228_r = node1220_r & pixel[126];
      node1228_l = node1220_r & ~pixel[126];
      node1229_r = node1228_l & pixel[623];
      node1229_l = node1228_l & ~pixel[623];
      node1230 = node1229_l;
      node1231 = node1229_r;
      node1232_r = node1228_r & pixel[430];
      node1232_l = node1228_r & ~pixel[430];
      node1233 = node1232_l;
      node1234 = node1232_r;
      node1235_r = node1203_r & pixel[126];
      node1235_l = node1203_r & ~pixel[126];
      node1236_r = node1235_l & pixel[156];
      node1236_l = node1235_l & ~pixel[156];
      node1237_r = node1236_l & pixel[684];
      node1237_l = node1236_l & ~pixel[684];
      node1238_r = node1237_l & pixel[96];
      node1238_l = node1237_l & ~pixel[96];
      node1239 = node1238_l;
      node1240 = node1238_r;
      node1241_r = node1237_r & pixel[218];
      node1241_l = node1237_r & ~pixel[218];
      node1242 = node1241_l;
      node1243 = node1241_r;
      node1244_r = node1236_r & pixel[656];
      node1244_l = node1236_r & ~pixel[656];
      node1245_r = node1244_l & pixel[100];
      node1245_l = node1244_l & ~pixel[100];
      node1246 = node1245_l;
      node1247 = node1245_r;
      node1248_r = node1244_r & pixel[455];
      node1248_l = node1244_r & ~pixel[455];
      node1249 = node1248_l;
      node1250 = node1248_r;
      node1251_r = node1235_r & pixel[659];
      node1251_l = node1235_r & ~pixel[659];
      node1252_r = node1251_l & pixel[236];
      node1252_l = node1251_l & ~pixel[236];
      node1253_r = node1252_l & pixel[495];
      node1253_l = node1252_l & ~pixel[495];
      node1254 = node1253_l;
      node1255 = node1253_r;
      node1256_r = node1252_r & pixel[662];
      node1256_l = node1252_r & ~pixel[662];
      node1257 = node1256_l;
      node1258 = node1256_r;
      node1259_r = node1251_r & pixel[400];
      node1259_l = node1251_r & ~pixel[400];
      node1260_r = node1259_l & pixel[580];
      node1260_l = node1259_l & ~pixel[580];
      node1261 = node1260_l;
      node1262 = node1260_r;
      node1263_r = node1259_r & pixel[211];
      node1263_l = node1259_r & ~pixel[211];
      node1264 = node1263_l;
      node1265 = node1263_r;
      node1266_r = node1202_r & pixel[624];
      node1266_l = node1202_r & ~pixel[624];
      node1267_r = node1266_l & pixel[153];
      node1267_l = node1266_l & ~pixel[153];
      node1268_r = node1267_l & pixel[238];
      node1268_l = node1267_l & ~pixel[238];
      node1269_r = node1268_l & pixel[340];
      node1269_l = node1268_l & ~pixel[340];
      node1270_r = node1269_l & pixel[266];
      node1270_l = node1269_l & ~pixel[266];
      node1271 = node1270_l;
      node1272 = node1270_r;
      node1273 = node1269_r;
      node1274_r = node1268_r & pixel[469];
      node1274_l = node1268_r & ~pixel[469];
      node1275_r = node1274_l & pixel[230];
      node1275_l = node1274_l & ~pixel[230];
      node1276 = node1275_l;
      node1277 = node1275_r;
      node1278_r = node1274_r & pixel[608];
      node1278_l = node1274_r & ~pixel[608];
      node1279 = node1278_l;
      node1280 = node1278_r;
      node1281_r = node1267_r & pixel[458];
      node1281_l = node1267_r & ~pixel[458];
      node1282_r = node1281_l & pixel[661];
      node1282_l = node1281_l & ~pixel[661];
      node1283_r = node1282_l & pixel[154];
      node1283_l = node1282_l & ~pixel[154];
      node1284 = node1283_l;
      node1285 = node1283_r;
      node1286_r = node1282_r & pixel[573];
      node1286_l = node1282_r & ~pixel[573];
      node1287 = node1286_l;
      node1288 = node1286_r;
      node1289_r = node1281_r & pixel[183];
      node1289_l = node1281_r & ~pixel[183];
      node1290_r = node1289_l & pixel[551];
      node1290_l = node1289_l & ~pixel[551];
      node1291 = node1290_l;
      node1292 = node1290_r;
      node1293_r = node1289_r & pixel[347];
      node1293_l = node1289_r & ~pixel[347];
      node1294 = node1293_l;
      node1295 = node1293_r;
      node1296_r = node1266_r & pixel[489];
      node1296_l = node1266_r & ~pixel[489];
      node1297_r = node1296_l & pixel[220];
      node1297_l = node1296_l & ~pixel[220];
      node1298_r = node1297_l & pixel[347];
      node1298_l = node1297_l & ~pixel[347];
      node1299_r = node1298_l & pixel[386];
      node1299_l = node1298_l & ~pixel[386];
      node1300 = node1299_l;
      node1301 = node1299_r;
      node1302_r = node1298_r & pixel[513];
      node1302_l = node1298_r & ~pixel[513];
      node1303 = node1302_l;
      node1304 = node1302_r;
      node1305_r = node1297_r & pixel[387];
      node1305_l = node1297_r & ~pixel[387];
      node1306_r = node1305_l & pixel[244];
      node1306_l = node1305_l & ~pixel[244];
      node1307 = node1306_l;
      node1308 = node1306_r;
      node1309 = node1305_r;
      node1310_r = node1296_r & pixel[713];
      node1310_l = node1296_r & ~pixel[713];
      node1311_r = node1310_l & pixel[263];
      node1311_l = node1310_l & ~pixel[263];
      node1312_r = node1311_l & pixel[464];
      node1312_l = node1311_l & ~pixel[464];
      node1313 = node1312_l;
      node1314 = node1312_r;
      node1315_r = node1311_r & pixel[539];
      node1315_l = node1311_r & ~pixel[539];
      node1316 = node1315_l;
      node1317 = node1315_r;
      node1318_r = node1310_r & pixel[321];
      node1318_l = node1310_r & ~pixel[321];
      node1319 = node1318_l;
      node1320 = node1318_r;
      node1321_r = node1201_r & pixel[513];
      node1321_l = node1201_r & ~pixel[513];
      node1322_r = node1321_l & pixel[386];
      node1322_l = node1321_l & ~pixel[386];
      node1323_r = node1322_l & pixel[353];
      node1323_l = node1322_l & ~pixel[353];
      node1324_r = node1323_l & pixel[190];
      node1324_l = node1323_l & ~pixel[190];
      node1325_r = node1324_l & pixel[217];
      node1325_l = node1324_l & ~pixel[217];
      node1326_r = node1325_l & pixel[150];
      node1326_l = node1325_l & ~pixel[150];
      node1327 = node1326_l;
      node1328 = node1326_r;
      node1329_r = node1325_r & pixel[481];
      node1329_l = node1325_r & ~pixel[481];
      node1330 = node1329_l;
      node1331 = node1329_r;
      node1332_r = node1324_r & pixel[413];
      node1332_l = node1324_r & ~pixel[413];
      node1333_r = node1332_l & pixel[205];
      node1333_l = node1332_l & ~pixel[205];
      node1334 = node1333_l;
      node1335 = node1333_r;
      node1336_r = node1332_r & pixel[639];
      node1336_l = node1332_r & ~pixel[639];
      node1337 = node1336_l;
      node1338 = node1336_r;
      node1339_r = node1323_r & pixel[375];
      node1339_l = node1323_r & ~pixel[375];
      node1340_r = node1339_l & pixel[483];
      node1340_l = node1339_l & ~pixel[483];
      node1341_r = node1340_l & pixel[712];
      node1341_l = node1340_l & ~pixel[712];
      node1342 = node1341_l;
      node1343 = node1341_r;
      node1344_r = node1340_r & pixel[152];
      node1344_l = node1340_r & ~pixel[152];
      node1345 = node1344_l;
      node1346 = node1344_r;
      node1347_r = node1339_r & pixel[272];
      node1347_l = node1339_r & ~pixel[272];
      node1348_r = node1347_l & pixel[174];
      node1348_l = node1347_l & ~pixel[174];
      node1349 = node1348_l;
      node1350 = node1348_r;
      node1351_r = node1347_r & pixel[207];
      node1351_l = node1347_r & ~pixel[207];
      node1352 = node1351_l;
      node1353 = node1351_r;
      node1354_r = node1322_r & pixel[382];
      node1354_l = node1322_r & ~pixel[382];
      node1355_r = node1354_l & pixel[635];
      node1355_l = node1354_l & ~pixel[635];
      node1356 = node1355_l;
      node1357_r = node1355_r & pixel[344];
      node1357_l = node1355_r & ~pixel[344];
      node1358_r = node1357_l & pixel[485];
      node1358_l = node1357_l & ~pixel[485];
      node1359 = node1358_l;
      node1360 = node1358_r;
      node1361 = node1357_r;
      node1362_r = node1354_r & pixel[202];
      node1362_l = node1354_r & ~pixel[202];
      node1363_r = node1362_l & pixel[373];
      node1363_l = node1362_l & ~pixel[373];
      node1364_r = node1363_l & pixel[499];
      node1364_l = node1363_l & ~pixel[499];
      node1365 = node1364_l;
      node1366 = node1364_r;
      node1367_r = node1363_r & pixel[321];
      node1367_l = node1363_r & ~pixel[321];
      node1368 = node1367_l;
      node1369 = node1367_r;
      node1370_r = node1362_r & pixel[540];
      node1370_l = node1362_r & ~pixel[540];
      node1371 = node1370_l;
      node1372 = node1370_r;
      node1373_r = node1321_r & pixel[274];
      node1373_l = node1321_r & ~pixel[274];
      node1374_r = node1373_l & pixel[299];
      node1374_l = node1373_l & ~pixel[299];
      node1375_r = node1374_l & pixel[486];
      node1375_l = node1374_l & ~pixel[486];
      node1376_r = node1375_l & pixel[624];
      node1376_l = node1375_l & ~pixel[624];
      node1377 = node1376_l;
      node1378_r = node1376_r & pixel[329];
      node1378_l = node1376_r & ~pixel[329];
      node1379 = node1378_l;
      node1380 = node1378_r;
      node1381_r = node1375_r & pixel[438];
      node1381_l = node1375_r & ~pixel[438];
      node1382_r = node1381_l & pixel[408];
      node1382_l = node1381_l & ~pixel[408];
      node1383 = node1382_l;
      node1384 = node1382_r;
      node1385_r = node1381_r & pixel[385];
      node1385_l = node1381_r & ~pixel[385];
      node1386 = node1385_l;
      node1387 = node1385_r;
      node1388_r = node1374_r & pixel[406];
      node1388_l = node1374_r & ~pixel[406];
      node1389_r = node1388_l & pixel[371];
      node1389_l = node1388_l & ~pixel[371];
      node1390 = node1389_l;
      node1391 = node1389_r;
      node1392_r = node1388_r & pixel[509];
      node1392_l = node1388_r & ~pixel[509];
      node1393_r = node1392_l & pixel[446];
      node1393_l = node1392_l & ~pixel[446];
      node1394 = node1393_l;
      node1395 = node1393_r;
      node1396 = node1392_r;
      node1397_r = node1373_r & pixel[413];
      node1397_l = node1373_r & ~pixel[413];
      node1398_r = node1397_l & pixel[372];
      node1398_l = node1397_l & ~pixel[372];
      node1399 = node1398_l;
      node1400_r = node1398_r & pixel[488];
      node1400_l = node1398_r & ~pixel[488];
      node1401_r = node1400_l & pixel[464];
      node1401_l = node1400_l & ~pixel[464];
      node1402 = node1401_l;
      node1403 = node1401_r;
      node1404_r = node1400_r & pixel[184];
      node1404_l = node1400_r & ~pixel[184];
      node1405 = node1404_l;
      node1406 = node1404_r;
      node1407_r = node1397_r & pixel[517];
      node1407_l = node1397_r & ~pixel[517];
      node1408_r = node1407_l & pixel[267];
      node1408_l = node1407_l & ~pixel[267];
      node1409 = node1408_l;
      node1410 = node1408_r;
      node1411_r = node1407_r & pixel[610];
      node1411_l = node1407_r & ~pixel[610];
      node1412_r = node1411_l & pixel[435];
      node1412_l = node1411_l & ~pixel[435];
      node1413 = node1412_l;
      node1414 = node1412_r;
      node1415 = node1411_r;
      node1416_r = node1200_r & pixel[656];
      node1416_l = node1200_r & ~pixel[656];
      node1417_r = node1416_l & pixel[189];
      node1417_l = node1416_l & ~pixel[189];
      node1418_r = node1417_l & pixel[269];
      node1418_l = node1417_l & ~pixel[269];
      node1419_r = node1418_l & pixel[243];
      node1419_l = node1418_l & ~pixel[243];
      node1420_r = node1419_l & pixel[609];
      node1420_l = node1419_l & ~pixel[609];
      node1421_r = node1420_l & pixel[458];
      node1421_l = node1420_l & ~pixel[458];
      node1422_r = node1421_l & pixel[355];
      node1422_l = node1421_l & ~pixel[355];
      node1423 = node1422_l;
      node1424 = node1422_r;
      node1425_r = node1421_r & pixel[247];
      node1425_l = node1421_r & ~pixel[247];
      node1426 = node1425_l;
      node1427 = node1425_r;
      node1428_r = node1420_r & pixel[173];
      node1428_l = node1420_r & ~pixel[173];
      node1429_r = node1428_l & pixel[344];
      node1429_l = node1428_l & ~pixel[344];
      node1430 = node1429_l;
      node1431 = node1429_r;
      node1432_r = node1428_r & pixel[597];
      node1432_l = node1428_r & ~pixel[597];
      node1433 = node1432_l;
      node1434 = node1432_r;
      node1435_r = node1419_r & pixel[679];
      node1435_l = node1419_r & ~pixel[679];
      node1436_r = node1435_l & pixel[596];
      node1436_l = node1435_l & ~pixel[596];
      node1437_r = node1436_l & pixel[320];
      node1437_l = node1436_l & ~pixel[320];
      node1438 = node1437_l;
      node1439 = node1437_r;
      node1440_r = node1436_r & pixel[275];
      node1440_l = node1436_r & ~pixel[275];
      node1441 = node1440_l;
      node1442 = node1440_r;
      node1443_r = node1435_r & pixel[459];
      node1443_l = node1435_r & ~pixel[459];
      node1444 = node1443_l;
      node1445_r = node1443_r & pixel[372];
      node1445_l = node1443_r & ~pixel[372];
      node1446 = node1445_l;
      node1447 = node1445_r;
      node1448_r = node1418_r & pixel[489];
      node1448_l = node1418_r & ~pixel[489];
      node1449_r = node1448_l & pixel[183];
      node1449_l = node1448_l & ~pixel[183];
      node1450_r = node1449_l & pixel[441];
      node1450_l = node1449_l & ~pixel[441];
      node1451_r = node1450_l & pixel[384];
      node1451_l = node1450_l & ~pixel[384];
      node1452 = node1451_l;
      node1453 = node1451_r;
      node1454_r = node1450_r & pixel[202];
      node1454_l = node1450_r & ~pixel[202];
      node1455 = node1454_l;
      node1456 = node1454_r;
      node1457_r = node1449_r & pixel[397];
      node1457_l = node1449_r & ~pixel[397];
      node1458_r = node1457_l & pixel[429];
      node1458_l = node1457_l & ~pixel[429];
      node1459 = node1458_l;
      node1460 = node1458_r;
      node1461_r = node1457_r & pixel[584];
      node1461_l = node1457_r & ~pixel[584];
      node1462 = node1461_l;
      node1463 = node1461_r;
      node1464_r = node1448_r & pixel[179];
      node1464_l = node1448_r & ~pixel[179];
      node1465_r = node1464_l & pixel[468];
      node1465_l = node1464_l & ~pixel[468];
      node1466_r = node1465_l & pixel[655];
      node1466_l = node1465_l & ~pixel[655];
      node1467 = node1466_l;
      node1468 = node1466_r;
      node1469_r = node1465_r & pixel[373];
      node1469_l = node1465_r & ~pixel[373];
      node1470 = node1469_l;
      node1471 = node1469_r;
      node1472_r = node1464_r & pixel[383];
      node1472_l = node1464_r & ~pixel[383];
      node1473_r = node1472_l & pixel[545];
      node1473_l = node1472_l & ~pixel[545];
      node1474 = node1473_l;
      node1475 = node1473_r;
      node1476_r = node1472_r & pixel[412];
      node1476_l = node1472_r & ~pixel[412];
      node1477 = node1476_l;
      node1478 = node1476_r;
      node1479_r = node1417_r & pixel[298];
      node1479_l = node1417_r & ~pixel[298];
      node1480_r = node1479_l & pixel[679];
      node1480_l = node1479_l & ~pixel[679];
      node1481_r = node1480_l & pixel[488];
      node1481_l = node1480_l & ~pixel[488];
      node1482_r = node1481_l & pixel[483];
      node1482_l = node1481_l & ~pixel[483];
      node1483_r = node1482_l & pixel[507];
      node1483_l = node1482_l & ~pixel[507];
      node1484 = node1483_l;
      node1485 = node1483_r;
      node1486_r = node1482_r & pixel[564];
      node1486_l = node1482_r & ~pixel[564];
      node1487 = node1486_l;
      node1488 = node1486_r;
      node1489_r = node1481_r & pixel[218];
      node1489_l = node1481_r & ~pixel[218];
      node1490_r = node1489_l & pixel[428];
      node1490_l = node1489_l & ~pixel[428];
      node1491 = node1490_l;
      node1492 = node1490_r;
      node1493_r = node1489_r & pixel[536];
      node1493_l = node1489_r & ~pixel[536];
      node1494 = node1493_l;
      node1495 = node1493_r;
      node1496_r = node1480_r & pixel[163];
      node1496_l = node1480_r & ~pixel[163];
      node1497_r = node1496_l & pixel[463];
      node1497_l = node1496_l & ~pixel[463];
      node1498 = node1497_l;
      node1499_r = node1497_r & pixel[204];
      node1499_l = node1497_r & ~pixel[204];
      node1500 = node1499_l;
      node1501 = node1499_r;
      node1502_r = node1496_r & pixel[510];
      node1502_l = node1496_r & ~pixel[510];
      node1503_r = node1502_l & pixel[521];
      node1503_l = node1502_l & ~pixel[521];
      node1504 = node1503_l;
      node1505 = node1503_r;
      node1506 = node1502_r;
      node1507_r = node1479_r & pixel[489];
      node1507_l = node1479_r & ~pixel[489];
      node1508_r = node1507_l & pixel[572];
      node1508_l = node1507_l & ~pixel[572];
      node1509 = node1508_l;
      node1510_r = node1508_r & pixel[427];
      node1510_l = node1508_r & ~pixel[427];
      node1511_r = node1510_l & pixel[485];
      node1511_l = node1510_l & ~pixel[485];
      node1512 = node1511_l;
      node1513 = node1511_r;
      node1514_r = node1510_r & pixel[235];
      node1514_l = node1510_r & ~pixel[235];
      node1515 = node1514_l;
      node1516 = node1514_r;
      node1517_r = node1507_r & pixel[211];
      node1517_l = node1507_r & ~pixel[211];
      node1518_r = node1517_l & pixel[357];
      node1518_l = node1517_l & ~pixel[357];
      node1519_r = node1518_l & pixel[537];
      node1519_l = node1518_l & ~pixel[537];
      node1520 = node1519_l;
      node1521 = node1519_r;
      node1522_r = node1518_r & pixel[510];
      node1522_l = node1518_r & ~pixel[510];
      node1523 = node1522_l;
      node1524 = node1522_r;
      node1525_r = node1517_r & pixel[595];
      node1525_l = node1517_r & ~pixel[595];
      node1526_r = node1525_l & pixel[300];
      node1526_l = node1525_l & ~pixel[300];
      node1527 = node1526_l;
      node1528 = node1526_r;
      node1529_r = node1525_r & pixel[580];
      node1529_l = node1525_r & ~pixel[580];
      node1530 = node1529_l;
      node1531 = node1529_r;
      node1532_r = node1416_r & pixel[439];
      node1532_l = node1416_r & ~pixel[439];
      node1533_r = node1532_l & pixel[325];
      node1533_l = node1532_l & ~pixel[325];
      node1534_r = node1533_l & pixel[462];
      node1534_l = node1533_l & ~pixel[462];
      node1535_r = node1534_l & pixel[385];
      node1535_l = node1534_l & ~pixel[385];
      node1536_r = node1535_l & pixel[460];
      node1536_l = node1535_l & ~pixel[460];
      node1537_r = node1536_l & pixel[152];
      node1537_l = node1536_l & ~pixel[152];
      node1538 = node1537_l;
      node1539 = node1537_r;
      node1540_r = node1536_r & pixel[217];
      node1540_l = node1536_r & ~pixel[217];
      node1541 = node1540_l;
      node1542 = node1540_r;
      node1543_r = node1535_r & pixel[271];
      node1543_l = node1535_r & ~pixel[271];
      node1544_r = node1543_l & pixel[354];
      node1544_l = node1543_l & ~pixel[354];
      node1545 = node1544_l;
      node1546 = node1544_r;
      node1547_r = node1543_r & pixel[689];
      node1547_l = node1543_r & ~pixel[689];
      node1548 = node1547_l;
      node1549 = node1547_r;
      node1550_r = node1534_r & pixel[383];
      node1550_l = node1534_r & ~pixel[383];
      node1551_r = node1550_l & pixel[191];
      node1551_l = node1550_l & ~pixel[191];
      node1552_r = node1551_l & pixel[293];
      node1552_l = node1551_l & ~pixel[293];
      node1553 = node1552_l;
      node1554 = node1552_r;
      node1555_r = node1551_r & pixel[381];
      node1555_l = node1551_r & ~pixel[381];
      node1556 = node1555_l;
      node1557 = node1555_r;
      node1558_r = node1550_r & pixel[735];
      node1558_l = node1550_r & ~pixel[735];
      node1559_r = node1558_l & pixel[710];
      node1559_l = node1558_l & ~pixel[710];
      node1560 = node1559_l;
      node1561 = node1559_r;
      node1562 = node1558_r;
      node1563_r = node1533_r & pixel[658];
      node1563_l = node1533_r & ~pixel[658];
      node1564_r = node1563_l & pixel[708];
      node1564_l = node1563_l & ~pixel[708];
      node1565_r = node1564_l & pixel[541];
      node1565_l = node1564_l & ~pixel[541];
      node1566_r = node1565_l & pixel[267];
      node1566_l = node1565_l & ~pixel[267];
      node1567 = node1566_l;
      node1568 = node1566_r;
      node1569_r = node1565_r & pixel[509];
      node1569_l = node1565_r & ~pixel[509];
      node1570 = node1569_l;
      node1571 = node1569_r;
      node1572_r = node1564_r & pixel[318];
      node1572_l = node1564_r & ~pixel[318];
      node1573_r = node1572_l & pixel[569];
      node1573_l = node1572_l & ~pixel[569];
      node1574 = node1573_l;
      node1575 = node1573_r;
      node1576_r = node1572_r & pixel[515];
      node1576_l = node1572_r & ~pixel[515];
      node1577 = node1576_l;
      node1578 = node1576_r;
      node1579_r = node1563_r & pixel[609];
      node1579_l = node1563_r & ~pixel[609];
      node1580_r = node1579_l & pixel[441];
      node1580_l = node1579_l & ~pixel[441];
      node1581_r = node1580_l & pixel[543];
      node1581_l = node1580_l & ~pixel[543];
      node1582 = node1581_l;
      node1583 = node1581_r;
      node1584_r = node1580_r & pixel[332];
      node1584_l = node1580_r & ~pixel[332];
      node1585 = node1584_l;
      node1586 = node1584_r;
      node1587_r = node1579_r & pixel[397];
      node1587_l = node1579_r & ~pixel[397];
      node1588_r = node1587_l & pixel[434];
      node1588_l = node1587_l & ~pixel[434];
      node1589 = node1588_l;
      node1590 = node1588_r;
      node1591 = node1587_r;
      node1592_r = node1532_r & pixel[462];
      node1592_l = node1532_r & ~pixel[462];
      node1593_r = node1592_l & pixel[296];
      node1593_l = node1592_l & ~pixel[296];
      node1594_r = node1593_l & pixel[515];
      node1594_l = node1593_l & ~pixel[515];
      node1595_r = node1594_l & pixel[456];
      node1595_l = node1594_l & ~pixel[456];
      node1596_r = node1595_l & pixel[295];
      node1596_l = node1595_l & ~pixel[295];
      node1597 = node1596_l;
      node1598 = node1596_r;
      node1599_r = node1595_r & pixel[383];
      node1599_l = node1595_r & ~pixel[383];
      node1600 = node1599_l;
      node1601 = node1599_r;
      node1602_r = node1594_r & pixel[380];
      node1602_l = node1594_r & ~pixel[380];
      node1603_r = node1602_l & pixel[244];
      node1603_l = node1602_l & ~pixel[244];
      node1604 = node1603_l;
      node1605 = node1603_r;
      node1606_r = node1602_r & pixel[599];
      node1606_l = node1602_r & ~pixel[599];
      node1607 = node1606_l;
      node1608 = node1606_r;
      node1609_r = node1593_r & pixel[484];
      node1609_l = node1593_r & ~pixel[484];
      node1610_r = node1609_l & pixel[653];
      node1610_l = node1609_l & ~pixel[653];
      node1611_r = node1610_l & pixel[459];
      node1611_l = node1610_l & ~pixel[459];
      node1612 = node1611_l;
      node1613 = node1611_r;
      node1614_r = node1610_r & pixel[263];
      node1614_l = node1610_r & ~pixel[263];
      node1615 = node1614_l;
      node1616 = node1614_r;
      node1617_r = node1609_r & pixel[301];
      node1617_l = node1609_r & ~pixel[301];
      node1618_r = node1617_l & pixel[401];
      node1618_l = node1617_l & ~pixel[401];
      node1619 = node1618_l;
      node1620 = node1618_r;
      node1621_r = node1617_r & pixel[330];
      node1621_l = node1617_r & ~pixel[330];
      node1622 = node1621_l;
      node1623 = node1621_r;
      node1624_r = node1592_r & pixel[659];
      node1624_l = node1592_r & ~pixel[659];
      node1625_r = node1624_l & pixel[330];
      node1625_l = node1624_l & ~pixel[330];
      node1626_r = node1625_l & pixel[184];
      node1626_l = node1625_l & ~pixel[184];
      node1627_r = node1626_l & pixel[576];
      node1627_l = node1626_l & ~pixel[576];
      node1628 = node1627_l;
      node1629 = node1627_r;
      node1630_r = node1626_r & pixel[522];
      node1630_l = node1626_r & ~pixel[522];
      node1631 = node1630_l;
      node1632 = node1630_r;
      node1633_r = node1625_r & pixel[156];
      node1633_l = node1625_r & ~pixel[156];
      node1634_r = node1633_l & pixel[432];
      node1634_l = node1633_l & ~pixel[432];
      node1635 = node1634_l;
      node1636 = node1634_r;
      node1637_r = node1633_r & pixel[186];
      node1637_l = node1633_r & ~pixel[186];
      node1638 = node1637_l;
      node1639 = node1637_r;
      node1640_r = node1624_r & pixel[593];
      node1640_l = node1624_r & ~pixel[593];
      node1641_r = node1640_l & pixel[487];
      node1641_l = node1640_l & ~pixel[487];
      node1642_r = node1641_l & pixel[330];
      node1642_l = node1641_l & ~pixel[330];
      node1643 = node1642_l;
      node1644 = node1642_r;
      node1645_r = node1641_r & pixel[182];
      node1645_l = node1641_r & ~pixel[182];
      node1646 = node1645_l;
      node1647 = node1645_r;
      node1648_r = node1640_r & pixel[687];
      node1648_l = node1640_r & ~pixel[687];
      node1649_r = node1648_l & pixel[541];
      node1649_l = node1648_l & ~pixel[541];
      node1650 = node1649_l;
      node1651 = node1649_r;
      node1652 = node1648_r;
      result0 = node14 | node42 | node58 | node60 | node75 | node78 | node108 | node122 | node130 | node134 | node135 | node138 | node150 | node151 | node154 | node158 | node168 | node184 | node197 | node216 | node343 | node347 | node368 | node369 | node380 | node384 | node387 | node388 | node397 | node400 | node403 | node404 | node406 | node424 | node430 | node451 | node468 | node488 | node500 | node501 | node505 | node507 | node508 | node513 | node515 | node592 | node634 | node645 | node646 | node662 | node668 | node672 | node676 | node677 | node689 | node701 | node709 | node711 | node713 | node721 | node722 | node724 | node725 | node729 | node747 | node835 | node839 | node1002 | node1132 | node1138 | node1163 | node1176 | node1309 | node1331 | node1356 | node1361 | node1369 | node1380 | node1390 | node1396 | node1402 | node1410 | node1413 | node1455 | node1462 | node1488 | node1515 | node1524 | node1545 | node1548 | node1586 | node1591 | node1605 | node1622 | node1623;
      result1 = node467 | node739 | node754 | node770 | node780 | node788 | node857 | node1223 | node1233 | node1258 | node1261;
      result2 = node18 | node49 | node83 | node86 | node102 | node103 | node112 | node119 | node141 | node163 | node182 | node190 | node193 | node196 | node199 | node200 | node206 | node211 | node233 | node235 | node247 | node248 | node262 | node281 | node292 | node307 | node308 | node313 | node321 | node324 | node326 | node329 | node342 | node344 | node353 | node355 | node366 | node381 | node407 | node427 | node433 | node446 | node455 | node463 | node476 | node477 | node520 | node521 | node533 | node536 | node537 | node544 | node552 | node553 | node555 | node556 | node559 | node570 | node572 | node582 | node586 | node589 | node609 | node610 | node614 | node617 | node649 | node652 | node663 | node666 | node691 | node715 | node758 | node764 | node765 | node777 | node781 | node795 | node806 | node818 | node826 | node829 | node841 | node845 | node849 | node864 | node867 | node886 | node900 | node915 | node922 | node930 | node931 | node934 | node937 | node944 | node945 | node947 | node952 | node959 | node969 | node975 | node978 | node979 | node983 | node986 | node1005 | node1009 | node1057 | node1067 | node1074 | node1078 | node1079 | node1093 | node1131 | node1144 | node1145 | node1155 | node1177 | node1183 | node1188 | node1189 | node1192 | node1196 | node1199 | node1239 | node1254 | node1366 | node1405 | node1415 | node1463 | node1470 | node1475 | node1477 | node1485 | node1495 | node1501 | node1531 | node1590 | node1629;
      result3 = node44 | node153 | node160 | node165 | node192 | node269 | node323 | node372 | node373 | node376 | node431 | node464 | node469 | node504 | node534 | node600 | node602 | node757 | node796 | node802 | node821 | node828 | node832 | node833 | node836 | node863 | node885 | node889 | node901 | node902 | node906 | node909 | node918 | node933 | node948 | node968 | node971 | node987 | node993 | node1003 | node1012 | node1028 | node1032 | node1035 | node1044 | node1047 | node1048 | node1056 | node1059 | node1066 | node1072 | node1075 | node1081 | node1089 | node1097 | node1099 | node1106 | node1118 | node1121 | node1122 | node1124 | node1133 | node1136 | node1148 | node1151 | node1152 | node1154 | node1160 | node1180 | node1181 | node1184 | node1191 | node1195 | node1198 | node1208 | node1216 | node1300 | node1303 | node1316 | node1328 | node1342 | node1345 | node1350 | node1353 | node1359 | node1371 | node1377 | node1391 | node1395 | node1433 | node1441 | node1453 | node1456 | node1459 | node1512 | node1589 | node1598 | node1612 | node1615 | node1616 | node1619 | node1632 | node1650;
      result4 = node11 | node21 | node26 | node68 | node89 | node93 | node98 | node101 | node111 | node126 | node174 | node212 | node215 | node225 | node226 | node229 | node243 | node261 | node274 | node276 | node311 | node328 | node356 | node418 | node434 | node445 | node483 | node523 | node527 | node540 | node541 | node577 | node621 | node648 | node655 | node700 | node716 | node742 | node750 | node785 | node805 | node810 | node813 | node817 | node822 | node846 | node870 | node877 | node1025 | node1026 | node1036 | node1040 | node1211 | node1224 | node1226 | node1234 | node1246 | node1250 | node1265 | node1271 | node1284 | node1291 | node1295 | node1427 | node1447 | node1520 | node1523 | node1527 | node1557 | node1567 | node1628 | node1631 | node1638;
      result5 = node17 | node29 | node32 | node45 | node55 | node67 | node74 | node120 | node157 | node161 | node167 | node208 | node228 | node236 | node241 | node250 | node258 | node266 | node268 | node337 | node351 | node365 | node375 | node383 | node390 | node396 | node399 | node414 | node415 | node480 | node487 | node490 | node498 | node563 | node583 | node599 | node603 | node615 | node630 | node671 | node675 | node743 | node746 | node749 | node755 | node771 | node789 | node879 | node888 | node892 | node905 | node908 | node956 | node960 | node1011 | node1018 | node1060 | node1063 | node1090 | node1092 | node1096 | node1100 | node1104 | node1109 | node1110 | node1113 | node1119 | node1127 | node1162 | node1167 | node1169 | node1175 | node1209 | node1215 | node1218 | node1219 | node1264 | node1308 | node1313 | node1320 | node1327 | node1330 | node1334 | node1335 | node1338 | node1343 | node1349 | node1352 | node1372 | node1379 | node1384 | node1386 | node1403 | node1423 | node1430 | node1442 | node1452 | node1467 | node1484 | node1487 | node1491 | node1494 | node1498 | node1505 | node1516 | node1521 | node1538 | node1539 | node1542 | node1546 | node1554 | node1556 | node1571 | node1585 | node1597 | node1600 | node1601 | node1604 | node1608 | node1643 | node1652;
      result6 = node20 | node28 | node36 | node41 | node52 | node61 | node71 | node77 | node92 | node99 | node107 | node110 | node127 | node129 | node137 | node142 | node144 | node145 | node175 | node177 | node178 | node189 | node204 | node207 | node217 | node232 | node240 | node252 | node259 | node277 | node283 | node284 | node297 | node312 | node320 | node330 | node335 | node346 | node352 | node391 | node421 | node440 | node442 | node443 | node450 | node454 | node461 | node473 | node484 | node497 | node510 | node514 | node528 | node543 | node585 | node590 | node607 | node618 | node622 | node624 | node625 | node631 | node633 | node638 | node656 | node688 | node693 | node702 | node705 | node706 | node726 | node740 | node778 | node803 | node812 | node842 | node848 | node984 | node999 | node1000 | node1006 | node1015 | node1016 | node1033 | node1043 | node1071 | node1240 | node1247 | node1255 | node1257 | node1292 | node1337 | node1424 | node1426 | node1431 | node1460 | node1471 | node1478 | node1492;
      result7 = node10 | node13 | node25 | node35 | node48 | node51 | node56 | node70 | node82 | node123 | node181 | node289 | node408 | node524 | node560 | node561 | node569 | node685 | node856 | node860 | node916 | node925 | node1272 | node1273 | node1277 | node1279 | node1562 | node1574 | node1635;
      result8 = node244 | node251 | node293 | node300 | node304 | node336 | node338 | node417 | node422 | node425 | node439 | node453 | node474 | node481 | node491 | node529 | node564 | node573 | node606 | node637 | node640 | node641 | node653 | node667 | node682 | node683 | node686 | node694 | node761 | node762 | node773 | node774 | node786 | node792 | node793 | node809 | node866 | node873 | node880 | node893 | node895 | node896 | node919 | node923 | node926 | node938 | node939 | node950 | node953 | node958 | node972 | node976 | node991 | node994 | node1019 | node1051 | node1064 | node1082 | node1112 | node1126 | node1137 | node1147 | node1159 | node1166 | node1170 | node1231 | node1243 | node1249 | node1262 | node1285 | node1287 | node1288 | node1304 | node1307 | node1314 | node1317 | node1346 | node1360 | node1365 | node1383 | node1387 | node1394 | node1399 | node1406 | node1409 | node1414 | node1434 | node1439 | node1474 | node1504 | node1506 | node1509 | node1513 | node1530 | node1541 | node1549 | node1553 | node1560 | node1561 | node1570 | node1575 | node1582 | node1583 | node1607 | node1613 | node1620 | node1639 | node1644 | node1646 | node1647 | node1651;
      result9 = node33 | node85 | node90 | node185 | node265 | node273 | node280 | node290 | node296 | node299 | node305 | node575 | node578 | node593 | node708 | node728 | node820 | node859 | node872 | node876 | node990 | node1029 | node1041 | node1050 | node1105 | node1212 | node1227 | node1230 | node1242 | node1276 | node1280 | node1294 | node1301 | node1319 | node1368 | node1438 | node1444 | node1446 | node1468 | node1500 | node1528 | node1568 | node1577 | node1578 | node1636;

      tree_3 = {result9, result8, result7, result6, result5, result4, result3, result2, result1, result0};
    end
  endfunction

  function [9:0] tree_4;
    input [783:0] pixel;

    reg node0_r;
    reg node0_l;
    reg node1_r;
    reg node1_l;
    reg node2_r;
    reg node2_l;
    reg node3_r;
    reg node3_l;
    reg node4_r;
    reg node4_l;
    reg node5_r;
    reg node5_l;
    reg node6_r;
    reg node6_l;
    reg node7_r;
    reg node7_l;
    reg node8_r;
    reg node8_l;
    reg node9_r;
    reg node9_l;
    reg node10;
    reg node11;
    reg node12_r;
    reg node12_l;
    reg node13;
    reg node14;
    reg node15_r;
    reg node15_l;
    reg node16_r;
    reg node16_l;
    reg node17;
    reg node18;
    reg node19_r;
    reg node19_l;
    reg node20;
    reg node21;
    reg node22_r;
    reg node22_l;
    reg node23;
    reg node24_r;
    reg node24_l;
    reg node25;
    reg node26;
    reg node27_r;
    reg node27_l;
    reg node28_r;
    reg node28_l;
    reg node29_r;
    reg node29_l;
    reg node30_r;
    reg node30_l;
    reg node31;
    reg node32;
    reg node33_r;
    reg node33_l;
    reg node34;
    reg node35;
    reg node36_r;
    reg node36_l;
    reg node37_r;
    reg node37_l;
    reg node38;
    reg node39;
    reg node40_r;
    reg node40_l;
    reg node41;
    reg node42;
    reg node43_r;
    reg node43_l;
    reg node44_r;
    reg node44_l;
    reg node45_r;
    reg node45_l;
    reg node46;
    reg node47;
    reg node48;
    reg node49;
    reg node50_r;
    reg node50_l;
    reg node51_r;
    reg node51_l;
    reg node52_r;
    reg node52_l;
    reg node53_r;
    reg node53_l;
    reg node54_r;
    reg node54_l;
    reg node55;
    reg node56;
    reg node57_r;
    reg node57_l;
    reg node58;
    reg node59;
    reg node60_r;
    reg node60_l;
    reg node61_r;
    reg node61_l;
    reg node62;
    reg node63;
    reg node64_r;
    reg node64_l;
    reg node65;
    reg node66;
    reg node67_r;
    reg node67_l;
    reg node68_r;
    reg node68_l;
    reg node69_r;
    reg node69_l;
    reg node70;
    reg node71;
    reg node72_r;
    reg node72_l;
    reg node73;
    reg node74;
    reg node75_r;
    reg node75_l;
    reg node76_r;
    reg node76_l;
    reg node77;
    reg node78;
    reg node79;
    reg node80_r;
    reg node80_l;
    reg node81_r;
    reg node81_l;
    reg node82_r;
    reg node82_l;
    reg node83_r;
    reg node83_l;
    reg node84;
    reg node85;
    reg node86_r;
    reg node86_l;
    reg node87;
    reg node88;
    reg node89_r;
    reg node89_l;
    reg node90_r;
    reg node90_l;
    reg node91;
    reg node92;
    reg node93_r;
    reg node93_l;
    reg node94;
    reg node95;
    reg node96_r;
    reg node96_l;
    reg node97_r;
    reg node97_l;
    reg node98_r;
    reg node98_l;
    reg node99;
    reg node100;
    reg node101_r;
    reg node101_l;
    reg node102;
    reg node103;
    reg node104_r;
    reg node104_l;
    reg node105_r;
    reg node105_l;
    reg node106;
    reg node107;
    reg node108_r;
    reg node108_l;
    reg node109;
    reg node110;
    reg node111_r;
    reg node111_l;
    reg node112_r;
    reg node112_l;
    reg node113_r;
    reg node113_l;
    reg node114_r;
    reg node114_l;
    reg node115_r;
    reg node115_l;
    reg node116_r;
    reg node116_l;
    reg node117;
    reg node118;
    reg node119_r;
    reg node119_l;
    reg node120;
    reg node121;
    reg node122_r;
    reg node122_l;
    reg node123_r;
    reg node123_l;
    reg node124;
    reg node125;
    reg node126_r;
    reg node126_l;
    reg node127;
    reg node128;
    reg node129_r;
    reg node129_l;
    reg node130_r;
    reg node130_l;
    reg node131_r;
    reg node131_l;
    reg node132;
    reg node133;
    reg node134_r;
    reg node134_l;
    reg node135;
    reg node136;
    reg node137_r;
    reg node137_l;
    reg node138_r;
    reg node138_l;
    reg node139;
    reg node140;
    reg node141_r;
    reg node141_l;
    reg node142;
    reg node143;
    reg node144_r;
    reg node144_l;
    reg node145_r;
    reg node145_l;
    reg node146_r;
    reg node146_l;
    reg node147_r;
    reg node147_l;
    reg node148;
    reg node149;
    reg node150_r;
    reg node150_l;
    reg node151;
    reg node152;
    reg node153_r;
    reg node153_l;
    reg node154_r;
    reg node154_l;
    reg node155;
    reg node156;
    reg node157_r;
    reg node157_l;
    reg node158;
    reg node159;
    reg node160_r;
    reg node160_l;
    reg node161_r;
    reg node161_l;
    reg node162_r;
    reg node162_l;
    reg node163;
    reg node164;
    reg node165_r;
    reg node165_l;
    reg node166;
    reg node167;
    reg node168_r;
    reg node168_l;
    reg node169_r;
    reg node169_l;
    reg node170;
    reg node171;
    reg node172_r;
    reg node172_l;
    reg node173;
    reg node174;
    reg node175_r;
    reg node175_l;
    reg node176_r;
    reg node176_l;
    reg node177_r;
    reg node177_l;
    reg node178_r;
    reg node178_l;
    reg node179_r;
    reg node179_l;
    reg node180;
    reg node181;
    reg node182_r;
    reg node182_l;
    reg node183;
    reg node184;
    reg node185_r;
    reg node185_l;
    reg node186_r;
    reg node186_l;
    reg node187;
    reg node188;
    reg node189_r;
    reg node189_l;
    reg node190;
    reg node191;
    reg node192_r;
    reg node192_l;
    reg node193_r;
    reg node193_l;
    reg node194;
    reg node195_r;
    reg node195_l;
    reg node196;
    reg node197;
    reg node198;
    reg node199;
    reg node200_r;
    reg node200_l;
    reg node201_r;
    reg node201_l;
    reg node202_r;
    reg node202_l;
    reg node203_r;
    reg node203_l;
    reg node204_r;
    reg node204_l;
    reg node205_r;
    reg node205_l;
    reg node206_r;
    reg node206_l;
    reg node207;
    reg node208;
    reg node209_r;
    reg node209_l;
    reg node210;
    reg node211;
    reg node212_r;
    reg node212_l;
    reg node213_r;
    reg node213_l;
    reg node214;
    reg node215;
    reg node216_r;
    reg node216_l;
    reg node217;
    reg node218;
    reg node219_r;
    reg node219_l;
    reg node220_r;
    reg node220_l;
    reg node221_r;
    reg node221_l;
    reg node222;
    reg node223;
    reg node224_r;
    reg node224_l;
    reg node225;
    reg node226;
    reg node227_r;
    reg node227_l;
    reg node228_r;
    reg node228_l;
    reg node229;
    reg node230;
    reg node231_r;
    reg node231_l;
    reg node232;
    reg node233;
    reg node234_r;
    reg node234_l;
    reg node235_r;
    reg node235_l;
    reg node236_r;
    reg node236_l;
    reg node237;
    reg node238_r;
    reg node238_l;
    reg node239;
    reg node240;
    reg node241_r;
    reg node241_l;
    reg node242;
    reg node243;
    reg node244_r;
    reg node244_l;
    reg node245_r;
    reg node245_l;
    reg node246;
    reg node247;
    reg node248;
    reg node249_r;
    reg node249_l;
    reg node250_r;
    reg node250_l;
    reg node251_r;
    reg node251_l;
    reg node252_r;
    reg node252_l;
    reg node253_r;
    reg node253_l;
    reg node254;
    reg node255;
    reg node256;
    reg node257_r;
    reg node257_l;
    reg node258;
    reg node259;
    reg node260_r;
    reg node260_l;
    reg node261_r;
    reg node261_l;
    reg node262_r;
    reg node262_l;
    reg node263;
    reg node264;
    reg node265;
    reg node266;
    reg node267_r;
    reg node267_l;
    reg node268;
    reg node269_r;
    reg node269_l;
    reg node270;
    reg node271;
    reg node272_r;
    reg node272_l;
    reg node273_r;
    reg node273_l;
    reg node274_r;
    reg node274_l;
    reg node275_r;
    reg node275_l;
    reg node276_r;
    reg node276_l;
    reg node277_r;
    reg node277_l;
    reg node278;
    reg node279;
    reg node280_r;
    reg node280_l;
    reg node281;
    reg node282;
    reg node283_r;
    reg node283_l;
    reg node284_r;
    reg node284_l;
    reg node285;
    reg node286;
    reg node287_r;
    reg node287_l;
    reg node288;
    reg node289;
    reg node290_r;
    reg node290_l;
    reg node291_r;
    reg node291_l;
    reg node292_r;
    reg node292_l;
    reg node293;
    reg node294;
    reg node295;
    reg node296_r;
    reg node296_l;
    reg node297_r;
    reg node297_l;
    reg node298;
    reg node299;
    reg node300_r;
    reg node300_l;
    reg node301;
    reg node302;
    reg node303_r;
    reg node303_l;
    reg node304_r;
    reg node304_l;
    reg node305_r;
    reg node305_l;
    reg node306;
    reg node307;
    reg node308_r;
    reg node308_l;
    reg node309_r;
    reg node309_l;
    reg node310;
    reg node311;
    reg node312_r;
    reg node312_l;
    reg node313;
    reg node314;
    reg node315_r;
    reg node315_l;
    reg node316_r;
    reg node316_l;
    reg node317_r;
    reg node317_l;
    reg node318;
    reg node319;
    reg node320_r;
    reg node320_l;
    reg node321;
    reg node322;
    reg node323_r;
    reg node323_l;
    reg node324_r;
    reg node324_l;
    reg node325;
    reg node326;
    reg node327_r;
    reg node327_l;
    reg node328;
    reg node329;
    reg node330_r;
    reg node330_l;
    reg node331_r;
    reg node331_l;
    reg node332_r;
    reg node332_l;
    reg node333_r;
    reg node333_l;
    reg node334_r;
    reg node334_l;
    reg node335;
    reg node336;
    reg node337;
    reg node338_r;
    reg node338_l;
    reg node339;
    reg node340;
    reg node341;
    reg node342_r;
    reg node342_l;
    reg node343_r;
    reg node343_l;
    reg node344_r;
    reg node344_l;
    reg node345_r;
    reg node345_l;
    reg node346;
    reg node347;
    reg node348;
    reg node349_r;
    reg node349_l;
    reg node350;
    reg node351_r;
    reg node351_l;
    reg node352;
    reg node353;
    reg node354_r;
    reg node354_l;
    reg node355;
    reg node356_r;
    reg node356_l;
    reg node357;
    reg node358;
    reg node359_r;
    reg node359_l;
    reg node360_r;
    reg node360_l;
    reg node361_r;
    reg node361_l;
    reg node362_r;
    reg node362_l;
    reg node363_r;
    reg node363_l;
    reg node364_r;
    reg node364_l;
    reg node365_r;
    reg node365_l;
    reg node366_r;
    reg node366_l;
    reg node367;
    reg node368;
    reg node369_r;
    reg node369_l;
    reg node370;
    reg node371;
    reg node372_r;
    reg node372_l;
    reg node373_r;
    reg node373_l;
    reg node374;
    reg node375;
    reg node376_r;
    reg node376_l;
    reg node377;
    reg node378;
    reg node379_r;
    reg node379_l;
    reg node380_r;
    reg node380_l;
    reg node381_r;
    reg node381_l;
    reg node382;
    reg node383;
    reg node384_r;
    reg node384_l;
    reg node385;
    reg node386;
    reg node387_r;
    reg node387_l;
    reg node388_r;
    reg node388_l;
    reg node389;
    reg node390;
    reg node391;
    reg node392_r;
    reg node392_l;
    reg node393_r;
    reg node393_l;
    reg node394_r;
    reg node394_l;
    reg node395_r;
    reg node395_l;
    reg node396;
    reg node397;
    reg node398_r;
    reg node398_l;
    reg node399;
    reg node400;
    reg node401_r;
    reg node401_l;
    reg node402_r;
    reg node402_l;
    reg node403;
    reg node404;
    reg node405_r;
    reg node405_l;
    reg node406;
    reg node407;
    reg node408_r;
    reg node408_l;
    reg node409_r;
    reg node409_l;
    reg node410_r;
    reg node410_l;
    reg node411;
    reg node412;
    reg node413_r;
    reg node413_l;
    reg node414;
    reg node415;
    reg node416_r;
    reg node416_l;
    reg node417;
    reg node418_r;
    reg node418_l;
    reg node419;
    reg node420;
    reg node421_r;
    reg node421_l;
    reg node422_r;
    reg node422_l;
    reg node423_r;
    reg node423_l;
    reg node424_r;
    reg node424_l;
    reg node425_r;
    reg node425_l;
    reg node426;
    reg node427;
    reg node428_r;
    reg node428_l;
    reg node429;
    reg node430;
    reg node431_r;
    reg node431_l;
    reg node432_r;
    reg node432_l;
    reg node433;
    reg node434;
    reg node435_r;
    reg node435_l;
    reg node436;
    reg node437;
    reg node438_r;
    reg node438_l;
    reg node439_r;
    reg node439_l;
    reg node440_r;
    reg node440_l;
    reg node441;
    reg node442;
    reg node443_r;
    reg node443_l;
    reg node444;
    reg node445;
    reg node446_r;
    reg node446_l;
    reg node447_r;
    reg node447_l;
    reg node448;
    reg node449;
    reg node450_r;
    reg node450_l;
    reg node451;
    reg node452;
    reg node453_r;
    reg node453_l;
    reg node454_r;
    reg node454_l;
    reg node455_r;
    reg node455_l;
    reg node456_r;
    reg node456_l;
    reg node457;
    reg node458;
    reg node459_r;
    reg node459_l;
    reg node460;
    reg node461;
    reg node462_r;
    reg node462_l;
    reg node463_r;
    reg node463_l;
    reg node464;
    reg node465;
    reg node466_r;
    reg node466_l;
    reg node467;
    reg node468;
    reg node469_r;
    reg node469_l;
    reg node470_r;
    reg node470_l;
    reg node471_r;
    reg node471_l;
    reg node472;
    reg node473;
    reg node474_r;
    reg node474_l;
    reg node475;
    reg node476;
    reg node477_r;
    reg node477_l;
    reg node478_r;
    reg node478_l;
    reg node479;
    reg node480;
    reg node481_r;
    reg node481_l;
    reg node482;
    reg node483;
    reg node484_r;
    reg node484_l;
    reg node485_r;
    reg node485_l;
    reg node486_r;
    reg node486_l;
    reg node487_r;
    reg node487_l;
    reg node488_r;
    reg node488_l;
    reg node489_r;
    reg node489_l;
    reg node490;
    reg node491;
    reg node492_r;
    reg node492_l;
    reg node493;
    reg node494;
    reg node495_r;
    reg node495_l;
    reg node496_r;
    reg node496_l;
    reg node497;
    reg node498;
    reg node499_r;
    reg node499_l;
    reg node500;
    reg node501;
    reg node502_r;
    reg node502_l;
    reg node503_r;
    reg node503_l;
    reg node504_r;
    reg node504_l;
    reg node505;
    reg node506;
    reg node507_r;
    reg node507_l;
    reg node508;
    reg node509;
    reg node510_r;
    reg node510_l;
    reg node511_r;
    reg node511_l;
    reg node512;
    reg node513;
    reg node514_r;
    reg node514_l;
    reg node515;
    reg node516;
    reg node517_r;
    reg node517_l;
    reg node518_r;
    reg node518_l;
    reg node519_r;
    reg node519_l;
    reg node520_r;
    reg node520_l;
    reg node521;
    reg node522;
    reg node523_r;
    reg node523_l;
    reg node524;
    reg node525;
    reg node526_r;
    reg node526_l;
    reg node527_r;
    reg node527_l;
    reg node528;
    reg node529;
    reg node530_r;
    reg node530_l;
    reg node531;
    reg node532;
    reg node533_r;
    reg node533_l;
    reg node534_r;
    reg node534_l;
    reg node535_r;
    reg node535_l;
    reg node536;
    reg node537;
    reg node538_r;
    reg node538_l;
    reg node539;
    reg node540;
    reg node541_r;
    reg node541_l;
    reg node542_r;
    reg node542_l;
    reg node543;
    reg node544;
    reg node545_r;
    reg node545_l;
    reg node546;
    reg node547;
    reg node548_r;
    reg node548_l;
    reg node549_r;
    reg node549_l;
    reg node550_r;
    reg node550_l;
    reg node551_r;
    reg node551_l;
    reg node552_r;
    reg node552_l;
    reg node553;
    reg node554;
    reg node555;
    reg node556_r;
    reg node556_l;
    reg node557;
    reg node558;
    reg node559_r;
    reg node559_l;
    reg node560_r;
    reg node560_l;
    reg node561;
    reg node562;
    reg node563;
    reg node564;
    reg node565_r;
    reg node565_l;
    reg node566_r;
    reg node566_l;
    reg node567_r;
    reg node567_l;
    reg node568_r;
    reg node568_l;
    reg node569_r;
    reg node569_l;
    reg node570_r;
    reg node570_l;
    reg node571_r;
    reg node571_l;
    reg node572;
    reg node573;
    reg node574_r;
    reg node574_l;
    reg node575;
    reg node576;
    reg node577_r;
    reg node577_l;
    reg node578_r;
    reg node578_l;
    reg node579;
    reg node580;
    reg node581_r;
    reg node581_l;
    reg node582;
    reg node583;
    reg node584_r;
    reg node584_l;
    reg node585_r;
    reg node585_l;
    reg node586_r;
    reg node586_l;
    reg node587;
    reg node588;
    reg node589_r;
    reg node589_l;
    reg node590;
    reg node591;
    reg node592_r;
    reg node592_l;
    reg node593_r;
    reg node593_l;
    reg node594;
    reg node595;
    reg node596_r;
    reg node596_l;
    reg node597;
    reg node598;
    reg node599_r;
    reg node599_l;
    reg node600_r;
    reg node600_l;
    reg node601_r;
    reg node601_l;
    reg node602_r;
    reg node602_l;
    reg node603;
    reg node604;
    reg node605_r;
    reg node605_l;
    reg node606;
    reg node607;
    reg node608_r;
    reg node608_l;
    reg node609_r;
    reg node609_l;
    reg node610;
    reg node611;
    reg node612_r;
    reg node612_l;
    reg node613;
    reg node614;
    reg node615_r;
    reg node615_l;
    reg node616_r;
    reg node616_l;
    reg node617_r;
    reg node617_l;
    reg node618;
    reg node619;
    reg node620_r;
    reg node620_l;
    reg node621;
    reg node622;
    reg node623_r;
    reg node623_l;
    reg node624_r;
    reg node624_l;
    reg node625;
    reg node626;
    reg node627_r;
    reg node627_l;
    reg node628;
    reg node629;
    reg node630_r;
    reg node630_l;
    reg node631_r;
    reg node631_l;
    reg node632_r;
    reg node632_l;
    reg node633_r;
    reg node633_l;
    reg node634_r;
    reg node634_l;
    reg node635;
    reg node636;
    reg node637_r;
    reg node637_l;
    reg node638;
    reg node639;
    reg node640_r;
    reg node640_l;
    reg node641_r;
    reg node641_l;
    reg node642;
    reg node643;
    reg node644_r;
    reg node644_l;
    reg node645;
    reg node646;
    reg node647_r;
    reg node647_l;
    reg node648_r;
    reg node648_l;
    reg node649_r;
    reg node649_l;
    reg node650;
    reg node651;
    reg node652_r;
    reg node652_l;
    reg node653;
    reg node654;
    reg node655_r;
    reg node655_l;
    reg node656_r;
    reg node656_l;
    reg node657;
    reg node658;
    reg node659_r;
    reg node659_l;
    reg node660;
    reg node661;
    reg node662_r;
    reg node662_l;
    reg node663_r;
    reg node663_l;
    reg node664_r;
    reg node664_l;
    reg node665_r;
    reg node665_l;
    reg node666;
    reg node667;
    reg node668_r;
    reg node668_l;
    reg node669;
    reg node670;
    reg node671_r;
    reg node671_l;
    reg node672_r;
    reg node672_l;
    reg node673;
    reg node674;
    reg node675_r;
    reg node675_l;
    reg node676;
    reg node677;
    reg node678_r;
    reg node678_l;
    reg node679_r;
    reg node679_l;
    reg node680;
    reg node681_r;
    reg node681_l;
    reg node682;
    reg node683;
    reg node684_r;
    reg node684_l;
    reg node685_r;
    reg node685_l;
    reg node686;
    reg node687;
    reg node688_r;
    reg node688_l;
    reg node689;
    reg node690;
    reg node691_r;
    reg node691_l;
    reg node692_r;
    reg node692_l;
    reg node693_r;
    reg node693_l;
    reg node694_r;
    reg node694_l;
    reg node695_r;
    reg node695_l;
    reg node696_r;
    reg node696_l;
    reg node697;
    reg node698;
    reg node699_r;
    reg node699_l;
    reg node700;
    reg node701;
    reg node702_r;
    reg node702_l;
    reg node703_r;
    reg node703_l;
    reg node704;
    reg node705;
    reg node706_r;
    reg node706_l;
    reg node707;
    reg node708;
    reg node709_r;
    reg node709_l;
    reg node710_r;
    reg node710_l;
    reg node711_r;
    reg node711_l;
    reg node712;
    reg node713;
    reg node714_r;
    reg node714_l;
    reg node715;
    reg node716;
    reg node717_r;
    reg node717_l;
    reg node718_r;
    reg node718_l;
    reg node719;
    reg node720;
    reg node721_r;
    reg node721_l;
    reg node722;
    reg node723;
    reg node724_r;
    reg node724_l;
    reg node725_r;
    reg node725_l;
    reg node726_r;
    reg node726_l;
    reg node727_r;
    reg node727_l;
    reg node728;
    reg node729;
    reg node730_r;
    reg node730_l;
    reg node731;
    reg node732;
    reg node733_r;
    reg node733_l;
    reg node734_r;
    reg node734_l;
    reg node735;
    reg node736;
    reg node737_r;
    reg node737_l;
    reg node738;
    reg node739;
    reg node740_r;
    reg node740_l;
    reg node741_r;
    reg node741_l;
    reg node742_r;
    reg node742_l;
    reg node743;
    reg node744;
    reg node745_r;
    reg node745_l;
    reg node746;
    reg node747;
    reg node748_r;
    reg node748_l;
    reg node749_r;
    reg node749_l;
    reg node750;
    reg node751;
    reg node752_r;
    reg node752_l;
    reg node753;
    reg node754;
    reg node755_r;
    reg node755_l;
    reg node756_r;
    reg node756_l;
    reg node757_r;
    reg node757_l;
    reg node758_r;
    reg node758_l;
    reg node759_r;
    reg node759_l;
    reg node760;
    reg node761;
    reg node762_r;
    reg node762_l;
    reg node763;
    reg node764;
    reg node765_r;
    reg node765_l;
    reg node766_r;
    reg node766_l;
    reg node767;
    reg node768;
    reg node769_r;
    reg node769_l;
    reg node770;
    reg node771;
    reg node772_r;
    reg node772_l;
    reg node773_r;
    reg node773_l;
    reg node774_r;
    reg node774_l;
    reg node775;
    reg node776;
    reg node777_r;
    reg node777_l;
    reg node778;
    reg node779;
    reg node780_r;
    reg node780_l;
    reg node781_r;
    reg node781_l;
    reg node782;
    reg node783;
    reg node784_r;
    reg node784_l;
    reg node785;
    reg node786;
    reg node787_r;
    reg node787_l;
    reg node788_r;
    reg node788_l;
    reg node789_r;
    reg node789_l;
    reg node790_r;
    reg node790_l;
    reg node791;
    reg node792;
    reg node793_r;
    reg node793_l;
    reg node794;
    reg node795;
    reg node796_r;
    reg node796_l;
    reg node797_r;
    reg node797_l;
    reg node798;
    reg node799;
    reg node800_r;
    reg node800_l;
    reg node801;
    reg node802;
    reg node803_r;
    reg node803_l;
    reg node804_r;
    reg node804_l;
    reg node805_r;
    reg node805_l;
    reg node806;
    reg node807;
    reg node808_r;
    reg node808_l;
    reg node809;
    reg node810;
    reg node811_r;
    reg node811_l;
    reg node812_r;
    reg node812_l;
    reg node813;
    reg node814;
    reg node815_r;
    reg node815_l;
    reg node816;
    reg node817;
    reg node818_r;
    reg node818_l;
    reg node819_r;
    reg node819_l;
    reg node820_r;
    reg node820_l;
    reg node821_r;
    reg node821_l;
    reg node822_r;
    reg node822_l;
    reg node823_r;
    reg node823_l;
    reg node824_r;
    reg node824_l;
    reg node825_r;
    reg node825_l;
    reg node826_r;
    reg node826_l;
    reg node827;
    reg node828;
    reg node829_r;
    reg node829_l;
    reg node830;
    reg node831;
    reg node832_r;
    reg node832_l;
    reg node833_r;
    reg node833_l;
    reg node834;
    reg node835;
    reg node836_r;
    reg node836_l;
    reg node837;
    reg node838;
    reg node839_r;
    reg node839_l;
    reg node840_r;
    reg node840_l;
    reg node841_r;
    reg node841_l;
    reg node842;
    reg node843;
    reg node844_r;
    reg node844_l;
    reg node845;
    reg node846;
    reg node847_r;
    reg node847_l;
    reg node848_r;
    reg node848_l;
    reg node849;
    reg node850;
    reg node851;
    reg node852_r;
    reg node852_l;
    reg node853_r;
    reg node853_l;
    reg node854_r;
    reg node854_l;
    reg node855_r;
    reg node855_l;
    reg node856;
    reg node857;
    reg node858_r;
    reg node858_l;
    reg node859;
    reg node860;
    reg node861_r;
    reg node861_l;
    reg node862_r;
    reg node862_l;
    reg node863;
    reg node864;
    reg node865_r;
    reg node865_l;
    reg node866;
    reg node867;
    reg node868_r;
    reg node868_l;
    reg node869_r;
    reg node869_l;
    reg node870_r;
    reg node870_l;
    reg node871;
    reg node872;
    reg node873;
    reg node874;
    reg node875_r;
    reg node875_l;
    reg node876_r;
    reg node876_l;
    reg node877_r;
    reg node877_l;
    reg node878_r;
    reg node878_l;
    reg node879_r;
    reg node879_l;
    reg node880;
    reg node881;
    reg node882_r;
    reg node882_l;
    reg node883;
    reg node884;
    reg node885_r;
    reg node885_l;
    reg node886_r;
    reg node886_l;
    reg node887;
    reg node888;
    reg node889_r;
    reg node889_l;
    reg node890;
    reg node891;
    reg node892_r;
    reg node892_l;
    reg node893_r;
    reg node893_l;
    reg node894_r;
    reg node894_l;
    reg node895;
    reg node896;
    reg node897_r;
    reg node897_l;
    reg node898;
    reg node899;
    reg node900_r;
    reg node900_l;
    reg node901_r;
    reg node901_l;
    reg node902;
    reg node903;
    reg node904_r;
    reg node904_l;
    reg node905;
    reg node906;
    reg node907_r;
    reg node907_l;
    reg node908_r;
    reg node908_l;
    reg node909_r;
    reg node909_l;
    reg node910_r;
    reg node910_l;
    reg node911;
    reg node912;
    reg node913_r;
    reg node913_l;
    reg node914;
    reg node915;
    reg node916_r;
    reg node916_l;
    reg node917_r;
    reg node917_l;
    reg node918;
    reg node919;
    reg node920_r;
    reg node920_l;
    reg node921;
    reg node922;
    reg node923_r;
    reg node923_l;
    reg node924_r;
    reg node924_l;
    reg node925_r;
    reg node925_l;
    reg node926;
    reg node927;
    reg node928_r;
    reg node928_l;
    reg node929;
    reg node930;
    reg node931_r;
    reg node931_l;
    reg node932_r;
    reg node932_l;
    reg node933;
    reg node934;
    reg node935_r;
    reg node935_l;
    reg node936;
    reg node937;
    reg node938_r;
    reg node938_l;
    reg node939_r;
    reg node939_l;
    reg node940_r;
    reg node940_l;
    reg node941_r;
    reg node941_l;
    reg node942_r;
    reg node942_l;
    reg node943_r;
    reg node943_l;
    reg node944;
    reg node945;
    reg node946_r;
    reg node946_l;
    reg node947;
    reg node948;
    reg node949_r;
    reg node949_l;
    reg node950;
    reg node951_r;
    reg node951_l;
    reg node952;
    reg node953;
    reg node954;
    reg node955_r;
    reg node955_l;
    reg node956_r;
    reg node956_l;
    reg node957_r;
    reg node957_l;
    reg node958;
    reg node959;
    reg node960_r;
    reg node960_l;
    reg node961;
    reg node962_r;
    reg node962_l;
    reg node963;
    reg node964;
    reg node965_r;
    reg node965_l;
    reg node966_r;
    reg node966_l;
    reg node967_r;
    reg node967_l;
    reg node968;
    reg node969;
    reg node970;
    reg node971;
    reg node972_r;
    reg node972_l;
    reg node973_r;
    reg node973_l;
    reg node974_r;
    reg node974_l;
    reg node975_r;
    reg node975_l;
    reg node976;
    reg node977_r;
    reg node977_l;
    reg node978;
    reg node979;
    reg node980_r;
    reg node980_l;
    reg node981_r;
    reg node981_l;
    reg node982;
    reg node983;
    reg node984;
    reg node985_r;
    reg node985_l;
    reg node986;
    reg node987;
    reg node988;
    reg node989_r;
    reg node989_l;
    reg node990_r;
    reg node990_l;
    reg node991_r;
    reg node991_l;
    reg node992_r;
    reg node992_l;
    reg node993_r;
    reg node993_l;
    reg node994_r;
    reg node994_l;
    reg node995_r;
    reg node995_l;
    reg node996;
    reg node997;
    reg node998_r;
    reg node998_l;
    reg node999;
    reg node1000;
    reg node1001_r;
    reg node1001_l;
    reg node1002_r;
    reg node1002_l;
    reg node1003;
    reg node1004;
    reg node1005_r;
    reg node1005_l;
    reg node1006;
    reg node1007;
    reg node1008_r;
    reg node1008_l;
    reg node1009_r;
    reg node1009_l;
    reg node1010_r;
    reg node1010_l;
    reg node1011;
    reg node1012;
    reg node1013_r;
    reg node1013_l;
    reg node1014;
    reg node1015;
    reg node1016_r;
    reg node1016_l;
    reg node1017_r;
    reg node1017_l;
    reg node1018;
    reg node1019;
    reg node1020_r;
    reg node1020_l;
    reg node1021;
    reg node1022;
    reg node1023_r;
    reg node1023_l;
    reg node1024_r;
    reg node1024_l;
    reg node1025_r;
    reg node1025_l;
    reg node1026_r;
    reg node1026_l;
    reg node1027;
    reg node1028;
    reg node1029_r;
    reg node1029_l;
    reg node1030;
    reg node1031;
    reg node1032_r;
    reg node1032_l;
    reg node1033_r;
    reg node1033_l;
    reg node1034;
    reg node1035;
    reg node1036;
    reg node1037;
    reg node1038_r;
    reg node1038_l;
    reg node1039_r;
    reg node1039_l;
    reg node1040_r;
    reg node1040_l;
    reg node1041_r;
    reg node1041_l;
    reg node1042_r;
    reg node1042_l;
    reg node1043;
    reg node1044;
    reg node1045_r;
    reg node1045_l;
    reg node1046;
    reg node1047;
    reg node1048;
    reg node1049_r;
    reg node1049_l;
    reg node1050_r;
    reg node1050_l;
    reg node1051;
    reg node1052_r;
    reg node1052_l;
    reg node1053;
    reg node1054;
    reg node1055_r;
    reg node1055_l;
    reg node1056;
    reg node1057;
    reg node1058_r;
    reg node1058_l;
    reg node1059_r;
    reg node1059_l;
    reg node1060_r;
    reg node1060_l;
    reg node1061;
    reg node1062;
    reg node1063_r;
    reg node1063_l;
    reg node1064_r;
    reg node1064_l;
    reg node1065;
    reg node1066;
    reg node1067;
    reg node1068_r;
    reg node1068_l;
    reg node1069;
    reg node1070_r;
    reg node1070_l;
    reg node1071;
    reg node1072_r;
    reg node1072_l;
    reg node1073;
    reg node1074;
    reg node1075_r;
    reg node1075_l;
    reg node1076_r;
    reg node1076_l;
    reg node1077_r;
    reg node1077_l;
    reg node1078_r;
    reg node1078_l;
    reg node1079_r;
    reg node1079_l;
    reg node1080_r;
    reg node1080_l;
    reg node1081;
    reg node1082;
    reg node1083;
    reg node1084_r;
    reg node1084_l;
    reg node1085_r;
    reg node1085_l;
    reg node1086;
    reg node1087;
    reg node1088_r;
    reg node1088_l;
    reg node1089;
    reg node1090;
    reg node1091_r;
    reg node1091_l;
    reg node1092_r;
    reg node1092_l;
    reg node1093_r;
    reg node1093_l;
    reg node1094;
    reg node1095;
    reg node1096_r;
    reg node1096_l;
    reg node1097;
    reg node1098;
    reg node1099_r;
    reg node1099_l;
    reg node1100_r;
    reg node1100_l;
    reg node1101;
    reg node1102;
    reg node1103;
    reg node1104_r;
    reg node1104_l;
    reg node1105_r;
    reg node1105_l;
    reg node1106_r;
    reg node1106_l;
    reg node1107_r;
    reg node1107_l;
    reg node1108;
    reg node1109;
    reg node1110_r;
    reg node1110_l;
    reg node1111;
    reg node1112;
    reg node1113_r;
    reg node1113_l;
    reg node1114_r;
    reg node1114_l;
    reg node1115;
    reg node1116;
    reg node1117_r;
    reg node1117_l;
    reg node1118;
    reg node1119;
    reg node1120_r;
    reg node1120_l;
    reg node1121_r;
    reg node1121_l;
    reg node1122_r;
    reg node1122_l;
    reg node1123;
    reg node1124;
    reg node1125_r;
    reg node1125_l;
    reg node1126;
    reg node1127;
    reg node1128_r;
    reg node1128_l;
    reg node1129_r;
    reg node1129_l;
    reg node1130;
    reg node1131;
    reg node1132_r;
    reg node1132_l;
    reg node1133;
    reg node1134;
    reg node1135_r;
    reg node1135_l;
    reg node1136_r;
    reg node1136_l;
    reg node1137_r;
    reg node1137_l;
    reg node1138_r;
    reg node1138_l;
    reg node1139_r;
    reg node1139_l;
    reg node1140;
    reg node1141;
    reg node1142_r;
    reg node1142_l;
    reg node1143;
    reg node1144;
    reg node1145_r;
    reg node1145_l;
    reg node1146;
    reg node1147_r;
    reg node1147_l;
    reg node1148;
    reg node1149;
    reg node1150_r;
    reg node1150_l;
    reg node1151_r;
    reg node1151_l;
    reg node1152_r;
    reg node1152_l;
    reg node1153;
    reg node1154;
    reg node1155;
    reg node1156_r;
    reg node1156_l;
    reg node1157_r;
    reg node1157_l;
    reg node1158;
    reg node1159;
    reg node1160_r;
    reg node1160_l;
    reg node1161;
    reg node1162;
    reg node1163_r;
    reg node1163_l;
    reg node1164_r;
    reg node1164_l;
    reg node1165;
    reg node1166;
    reg node1167_r;
    reg node1167_l;
    reg node1168_r;
    reg node1168_l;
    reg node1169_r;
    reg node1169_l;
    reg node1170;
    reg node1171;
    reg node1172;
    reg node1173;
    reg node1174_r;
    reg node1174_l;
    reg node1175_r;
    reg node1175_l;
    reg node1176_r;
    reg node1176_l;
    reg node1177_r;
    reg node1177_l;
    reg node1178_r;
    reg node1178_l;
    reg node1179_r;
    reg node1179_l;
    reg node1180_r;
    reg node1180_l;
    reg node1181_r;
    reg node1181_l;
    reg node1182;
    reg node1183;
    reg node1184_r;
    reg node1184_l;
    reg node1185;
    reg node1186;
    reg node1187_r;
    reg node1187_l;
    reg node1188_r;
    reg node1188_l;
    reg node1189;
    reg node1190;
    reg node1191_r;
    reg node1191_l;
    reg node1192;
    reg node1193;
    reg node1194_r;
    reg node1194_l;
    reg node1195_r;
    reg node1195_l;
    reg node1196_r;
    reg node1196_l;
    reg node1197;
    reg node1198;
    reg node1199;
    reg node1200;
    reg node1201_r;
    reg node1201_l;
    reg node1202_r;
    reg node1202_l;
    reg node1203_r;
    reg node1203_l;
    reg node1204_r;
    reg node1204_l;
    reg node1205;
    reg node1206;
    reg node1207_r;
    reg node1207_l;
    reg node1208;
    reg node1209;
    reg node1210_r;
    reg node1210_l;
    reg node1211_r;
    reg node1211_l;
    reg node1212;
    reg node1213;
    reg node1214_r;
    reg node1214_l;
    reg node1215;
    reg node1216;
    reg node1217_r;
    reg node1217_l;
    reg node1218_r;
    reg node1218_l;
    reg node1219_r;
    reg node1219_l;
    reg node1220;
    reg node1221;
    reg node1222_r;
    reg node1222_l;
    reg node1223;
    reg node1224;
    reg node1225_r;
    reg node1225_l;
    reg node1226_r;
    reg node1226_l;
    reg node1227;
    reg node1228;
    reg node1229_r;
    reg node1229_l;
    reg node1230;
    reg node1231;
    reg node1232_r;
    reg node1232_l;
    reg node1233_r;
    reg node1233_l;
    reg node1234_r;
    reg node1234_l;
    reg node1235_r;
    reg node1235_l;
    reg node1236_r;
    reg node1236_l;
    reg node1237;
    reg node1238;
    reg node1239_r;
    reg node1239_l;
    reg node1240;
    reg node1241;
    reg node1242_r;
    reg node1242_l;
    reg node1243_r;
    reg node1243_l;
    reg node1244;
    reg node1245;
    reg node1246_r;
    reg node1246_l;
    reg node1247;
    reg node1248;
    reg node1249_r;
    reg node1249_l;
    reg node1250_r;
    reg node1250_l;
    reg node1251_r;
    reg node1251_l;
    reg node1252;
    reg node1253;
    reg node1254_r;
    reg node1254_l;
    reg node1255;
    reg node1256;
    reg node1257_r;
    reg node1257_l;
    reg node1258_r;
    reg node1258_l;
    reg node1259;
    reg node1260;
    reg node1261_r;
    reg node1261_l;
    reg node1262;
    reg node1263;
    reg node1264_r;
    reg node1264_l;
    reg node1265_r;
    reg node1265_l;
    reg node1266_r;
    reg node1266_l;
    reg node1267_r;
    reg node1267_l;
    reg node1268;
    reg node1269;
    reg node1270_r;
    reg node1270_l;
    reg node1271;
    reg node1272;
    reg node1273_r;
    reg node1273_l;
    reg node1274_r;
    reg node1274_l;
    reg node1275;
    reg node1276;
    reg node1277_r;
    reg node1277_l;
    reg node1278;
    reg node1279;
    reg node1280_r;
    reg node1280_l;
    reg node1281_r;
    reg node1281_l;
    reg node1282_r;
    reg node1282_l;
    reg node1283;
    reg node1284;
    reg node1285_r;
    reg node1285_l;
    reg node1286;
    reg node1287;
    reg node1288_r;
    reg node1288_l;
    reg node1289_r;
    reg node1289_l;
    reg node1290;
    reg node1291;
    reg node1292_r;
    reg node1292_l;
    reg node1293;
    reg node1294;
    reg node1295_r;
    reg node1295_l;
    reg node1296_r;
    reg node1296_l;
    reg node1297_r;
    reg node1297_l;
    reg node1298_r;
    reg node1298_l;
    reg node1299_r;
    reg node1299_l;
    reg node1300_r;
    reg node1300_l;
    reg node1301;
    reg node1302;
    reg node1303_r;
    reg node1303_l;
    reg node1304;
    reg node1305;
    reg node1306_r;
    reg node1306_l;
    reg node1307_r;
    reg node1307_l;
    reg node1308;
    reg node1309;
    reg node1310_r;
    reg node1310_l;
    reg node1311;
    reg node1312;
    reg node1313_r;
    reg node1313_l;
    reg node1314_r;
    reg node1314_l;
    reg node1315_r;
    reg node1315_l;
    reg node1316;
    reg node1317;
    reg node1318_r;
    reg node1318_l;
    reg node1319;
    reg node1320;
    reg node1321_r;
    reg node1321_l;
    reg node1322_r;
    reg node1322_l;
    reg node1323;
    reg node1324;
    reg node1325;
    reg node1326_r;
    reg node1326_l;
    reg node1327_r;
    reg node1327_l;
    reg node1328_r;
    reg node1328_l;
    reg node1329_r;
    reg node1329_l;
    reg node1330;
    reg node1331;
    reg node1332_r;
    reg node1332_l;
    reg node1333;
    reg node1334;
    reg node1335_r;
    reg node1335_l;
    reg node1336_r;
    reg node1336_l;
    reg node1337;
    reg node1338;
    reg node1339_r;
    reg node1339_l;
    reg node1340;
    reg node1341;
    reg node1342_r;
    reg node1342_l;
    reg node1343_r;
    reg node1343_l;
    reg node1344_r;
    reg node1344_l;
    reg node1345;
    reg node1346;
    reg node1347_r;
    reg node1347_l;
    reg node1348;
    reg node1349;
    reg node1350_r;
    reg node1350_l;
    reg node1351_r;
    reg node1351_l;
    reg node1352;
    reg node1353;
    reg node1354_r;
    reg node1354_l;
    reg node1355;
    reg node1356;
    reg node1357_r;
    reg node1357_l;
    reg node1358_r;
    reg node1358_l;
    reg node1359_r;
    reg node1359_l;
    reg node1360_r;
    reg node1360_l;
    reg node1361_r;
    reg node1361_l;
    reg node1362;
    reg node1363;
    reg node1364_r;
    reg node1364_l;
    reg node1365;
    reg node1366;
    reg node1367;
    reg node1368_r;
    reg node1368_l;
    reg node1369_r;
    reg node1369_l;
    reg node1370_r;
    reg node1370_l;
    reg node1371;
    reg node1372;
    reg node1373_r;
    reg node1373_l;
    reg node1374;
    reg node1375;
    reg node1376_r;
    reg node1376_l;
    reg node1377_r;
    reg node1377_l;
    reg node1378;
    reg node1379;
    reg node1380_r;
    reg node1380_l;
    reg node1381;
    reg node1382;
    reg node1383_r;
    reg node1383_l;
    reg node1384_r;
    reg node1384_l;
    reg node1385_r;
    reg node1385_l;
    reg node1386_r;
    reg node1386_l;
    reg node1387;
    reg node1388;
    reg node1389_r;
    reg node1389_l;
    reg node1390;
    reg node1391;
    reg node1392_r;
    reg node1392_l;
    reg node1393_r;
    reg node1393_l;
    reg node1394;
    reg node1395;
    reg node1396_r;
    reg node1396_l;
    reg node1397;
    reg node1398;
    reg node1399_r;
    reg node1399_l;
    reg node1400_r;
    reg node1400_l;
    reg node1401_r;
    reg node1401_l;
    reg node1402;
    reg node1403;
    reg node1404_r;
    reg node1404_l;
    reg node1405;
    reg node1406;
    reg node1407_r;
    reg node1407_l;
    reg node1408_r;
    reg node1408_l;
    reg node1409;
    reg node1410;
    reg node1411_r;
    reg node1411_l;
    reg node1412;
    reg node1413;
    reg node1414_r;
    reg node1414_l;
    reg node1415_r;
    reg node1415_l;
    reg node1416_r;
    reg node1416_l;
    reg node1417_r;
    reg node1417_l;
    reg node1418_r;
    reg node1418_l;
    reg node1419_r;
    reg node1419_l;
    reg node1420_r;
    reg node1420_l;
    reg node1421;
    reg node1422;
    reg node1423_r;
    reg node1423_l;
    reg node1424;
    reg node1425;
    reg node1426;
    reg node1427_r;
    reg node1427_l;
    reg node1428_r;
    reg node1428_l;
    reg node1429_r;
    reg node1429_l;
    reg node1430;
    reg node1431;
    reg node1432;
    reg node1433_r;
    reg node1433_l;
    reg node1434_r;
    reg node1434_l;
    reg node1435;
    reg node1436;
    reg node1437_r;
    reg node1437_l;
    reg node1438;
    reg node1439;
    reg node1440_r;
    reg node1440_l;
    reg node1441;
    reg node1442;
    reg node1443_r;
    reg node1443_l;
    reg node1444_r;
    reg node1444_l;
    reg node1445_r;
    reg node1445_l;
    reg node1446;
    reg node1447;
    reg node1448_r;
    reg node1448_l;
    reg node1449_r;
    reg node1449_l;
    reg node1450_r;
    reg node1450_l;
    reg node1451;
    reg node1452;
    reg node1453;
    reg node1454_r;
    reg node1454_l;
    reg node1455;
    reg node1456;
    reg node1457_r;
    reg node1457_l;
    reg node1458_r;
    reg node1458_l;
    reg node1459_r;
    reg node1459_l;
    reg node1460;
    reg node1461;
    reg node1462;
    reg node1463_r;
    reg node1463_l;
    reg node1464_r;
    reg node1464_l;
    reg node1465;
    reg node1466;
    reg node1467;
    reg node1468_r;
    reg node1468_l;
    reg node1469_r;
    reg node1469_l;
    reg node1470_r;
    reg node1470_l;
    reg node1471_r;
    reg node1471_l;
    reg node1472_r;
    reg node1472_l;
    reg node1473_r;
    reg node1473_l;
    reg node1474;
    reg node1475;
    reg node1476_r;
    reg node1476_l;
    reg node1477;
    reg node1478;
    reg node1479_r;
    reg node1479_l;
    reg node1480_r;
    reg node1480_l;
    reg node1481;
    reg node1482;
    reg node1483;
    reg node1484_r;
    reg node1484_l;
    reg node1485;
    reg node1486;
    reg node1487_r;
    reg node1487_l;
    reg node1488_r;
    reg node1488_l;
    reg node1489_r;
    reg node1489_l;
    reg node1490_r;
    reg node1490_l;
    reg node1491;
    reg node1492;
    reg node1493;
    reg node1494_r;
    reg node1494_l;
    reg node1495;
    reg node1496_r;
    reg node1496_l;
    reg node1497;
    reg node1498;
    reg node1499;
    reg node1500_r;
    reg node1500_l;
    reg node1501_r;
    reg node1501_l;
    reg node1502_r;
    reg node1502_l;
    reg node1503;
    reg node1504;
    reg node1505_r;
    reg node1505_l;
    reg node1506;
    reg node1507_r;
    reg node1507_l;
    reg node1508_r;
    reg node1508_l;
    reg node1509;
    reg node1510;
    reg node1511;
    reg node1512_r;
    reg node1512_l;
    reg node1513_r;
    reg node1513_l;
    reg node1514;
    reg node1515;
    reg node1516_r;
    reg node1516_l;
    reg node1517;
    reg node1518_r;
    reg node1518_l;
    reg node1519_r;
    reg node1519_l;
    reg node1520;
    reg node1521;
    reg node1522;
    reg result0;
    reg result1;
    reg result2;
    reg result3;
    reg result4;
    reg result5;
    reg result6;
    reg result7;
    reg result8;
    reg result9;

    begin
      node0_r = pixel[539];
      node0_l = ~pixel[539];
      node1_r = node0_l & pixel[433];
      node1_l = node0_l & ~pixel[433];
      node2_r = node1_l & pixel[257];
      node2_l = node1_l & ~pixel[257];
      node3_r = node2_l & pixel[376];
      node3_l = node2_l & ~pixel[376];
      node4_r = node3_l & pixel[181];
      node4_l = node3_l & ~pixel[181];
      node5_r = node4_l & pixel[238];
      node5_l = node4_l & ~pixel[238];
      node6_r = node5_l & pixel[68];
      node6_l = node5_l & ~pixel[68];
      node7_r = node6_l & pixel[293];
      node7_l = node6_l & ~pixel[293];
      node8_r = node7_l & pixel[574];
      node8_l = node7_l & ~pixel[574];
      node9_r = node8_l & pixel[567];
      node9_l = node8_l & ~pixel[567];
      node10 = node9_l;
      node11 = node9_r;
      node12_r = node8_r & pixel[414];
      node12_l = node8_r & ~pixel[414];
      node13 = node12_l;
      node14 = node12_r;
      node15_r = node7_r & pixel[290];
      node15_l = node7_r & ~pixel[290];
      node16_r = node15_l & pixel[129];
      node16_l = node15_l & ~pixel[129];
      node17 = node16_l;
      node18 = node16_r;
      node19_r = node15_r & pixel[512];
      node19_l = node15_r & ~pixel[512];
      node20 = node19_l;
      node21 = node19_r;
      node22_r = node6_r & pixel[155];
      node22_l = node6_r & ~pixel[155];
      node23 = node22_l;
      node24_r = node22_r & pixel[205];
      node24_l = node22_r & ~pixel[205];
      node25 = node24_l;
      node26 = node24_r;
      node27_r = node5_r & pixel[564];
      node27_l = node5_r & ~pixel[564];
      node28_r = node27_l & pixel[409];
      node28_l = node27_l & ~pixel[409];
      node29_r = node28_l & pixel[402];
      node29_l = node28_l & ~pixel[402];
      node30_r = node29_l & pixel[470];
      node30_l = node29_l & ~pixel[470];
      node31 = node30_l;
      node32 = node30_r;
      node33_r = node29_r & pixel[356];
      node33_l = node29_r & ~pixel[356];
      node34 = node33_l;
      node35 = node33_r;
      node36_r = node28_r & pixel[578];
      node36_l = node28_r & ~pixel[578];
      node37_r = node36_l & pixel[541];
      node37_l = node36_l & ~pixel[541];
      node38 = node37_l;
      node39 = node37_r;
      node40_r = node36_r & pixel[487];
      node40_l = node36_r & ~pixel[487];
      node41 = node40_l;
      node42 = node40_r;
      node43_r = node27_r & pixel[372];
      node43_l = node27_r & ~pixel[372];
      node44_r = node43_l & pixel[457];
      node44_l = node43_l & ~pixel[457];
      node45_r = node44_l & pixel[262];
      node45_l = node44_l & ~pixel[262];
      node46 = node45_l;
      node47 = node45_r;
      node48 = node44_r;
      node49 = node43_r;
      node50_r = node4_r & pixel[153];
      node50_l = node4_r & ~pixel[153];
      node51_r = node50_l & pixel[429];
      node51_l = node50_l & ~pixel[429];
      node52_r = node51_l & pixel[565];
      node52_l = node51_l & ~pixel[565];
      node53_r = node52_l & pixel[577];
      node53_l = node52_l & ~pixel[577];
      node54_r = node53_l & pixel[468];
      node54_l = node53_l & ~pixel[468];
      node55 = node54_l;
      node56 = node54_r;
      node57_r = node53_r & pixel[297];
      node57_l = node53_r & ~pixel[297];
      node58 = node57_l;
      node59 = node57_r;
      node60_r = node52_r & pixel[350];
      node60_l = node52_r & ~pixel[350];
      node61_r = node60_l & pixel[205];
      node61_l = node60_l & ~pixel[205];
      node62 = node61_l;
      node63 = node61_r;
      node64_r = node60_r & pixel[713];
      node64_l = node60_r & ~pixel[713];
      node65 = node64_l;
      node66 = node64_r;
      node67_r = node51_r & pixel[409];
      node67_l = node51_r & ~pixel[409];
      node68_r = node67_l & pixel[569];
      node68_l = node67_l & ~pixel[569];
      node69_r = node68_l & pixel[357];
      node69_l = node68_l & ~pixel[357];
      node70 = node69_l;
      node71 = node69_r;
      node72_r = node68_r & pixel[464];
      node72_l = node68_r & ~pixel[464];
      node73 = node72_l;
      node74 = node72_r;
      node75_r = node67_r & pixel[99];
      node75_l = node67_r & ~pixel[99];
      node76_r = node75_l & pixel[191];
      node76_l = node75_l & ~pixel[191];
      node77 = node76_l;
      node78 = node76_r;
      node79 = node75_r;
      node80_r = node50_r & pixel[242];
      node80_l = node50_r & ~pixel[242];
      node81_r = node80_l & pixel[519];
      node81_l = node80_l & ~pixel[519];
      node82_r = node81_l & pixel[463];
      node82_l = node81_l & ~pixel[463];
      node83_r = node82_l & pixel[458];
      node83_l = node82_l & ~pixel[458];
      node84 = node83_l;
      node85 = node83_r;
      node86_r = node82_r & pixel[290];
      node86_l = node82_r & ~pixel[290];
      node87 = node86_l;
      node88 = node86_r;
      node89_r = node81_r & pixel[545];
      node89_l = node81_r & ~pixel[545];
      node90_r = node89_l & pixel[401];
      node90_l = node89_l & ~pixel[401];
      node91 = node90_l;
      node92 = node90_r;
      node93_r = node89_r & pixel[627];
      node93_l = node89_r & ~pixel[627];
      node94 = node93_l;
      node95 = node93_r;
      node96_r = node80_r & pixel[491];
      node96_l = node80_r & ~pixel[491];
      node97_r = node96_l & pixel[512];
      node97_l = node96_l & ~pixel[512];
      node98_r = node97_l & pixel[295];
      node98_l = node97_l & ~pixel[295];
      node99 = node98_l;
      node100 = node98_r;
      node101_r = node97_r & pixel[488];
      node101_l = node97_r & ~pixel[488];
      node102 = node101_l;
      node103 = node101_r;
      node104_r = node96_r & pixel[572];
      node104_l = node96_r & ~pixel[572];
      node105_r = node104_l & pixel[327];
      node105_l = node104_l & ~pixel[327];
      node106 = node105_l;
      node107 = node105_r;
      node108_r = node104_r & pixel[399];
      node108_l = node104_r & ~pixel[399];
      node109 = node108_l;
      node110 = node108_r;
      node111_r = node3_r & pixel[101];
      node111_l = node3_r & ~pixel[101];
      node112_r = node111_l & pixel[296];
      node112_l = node111_l & ~pixel[296];
      node113_r = node112_l & pixel[458];
      node113_l = node112_l & ~pixel[458];
      node114_r = node113_l & pixel[517];
      node114_l = node113_l & ~pixel[517];
      node115_r = node114_l & pixel[297];
      node115_l = node114_l & ~pixel[297];
      node116_r = node115_l & pixel[267];
      node116_l = node115_l & ~pixel[267];
      node117 = node116_l;
      node118 = node116_r;
      node119_r = node115_r & pixel[624];
      node119_l = node115_r & ~pixel[624];
      node120 = node119_l;
      node121 = node119_r;
      node122_r = node114_r & pixel[326];
      node122_l = node114_r & ~pixel[326];
      node123_r = node122_l & pixel[377];
      node123_l = node122_l & ~pixel[377];
      node124 = node123_l;
      node125 = node123_r;
      node126_r = node122_r & pixel[522];
      node126_l = node122_r & ~pixel[522];
      node127 = node126_l;
      node128 = node126_r;
      node129_r = node113_r & pixel[300];
      node129_l = node113_r & ~pixel[300];
      node130_r = node129_l & pixel[297];
      node130_l = node129_l & ~pixel[297];
      node131_r = node130_l & pixel[544];
      node131_l = node130_l & ~pixel[544];
      node132 = node131_l;
      node133 = node131_r;
      node134_r = node130_r & pixel[598];
      node134_l = node130_r & ~pixel[598];
      node135 = node134_l;
      node136 = node134_r;
      node137_r = node129_r & pixel[351];
      node137_l = node129_r & ~pixel[351];
      node138_r = node137_l & pixel[186];
      node138_l = node137_l & ~pixel[186];
      node139 = node138_l;
      node140 = node138_r;
      node141_r = node137_r & pixel[372];
      node141_l = node137_r & ~pixel[372];
      node142 = node141_l;
      node143 = node141_r;
      node144_r = node112_r & pixel[180];
      node144_l = node112_r & ~pixel[180];
      node145_r = node144_l & pixel[273];
      node145_l = node144_l & ~pixel[273];
      node146_r = node145_l & pixel[459];
      node146_l = node145_l & ~pixel[459];
      node147_r = node146_l & pixel[155];
      node147_l = node146_l & ~pixel[155];
      node148 = node147_l;
      node149 = node147_r;
      node150_r = node146_r & pixel[191];
      node150_l = node146_r & ~pixel[191];
      node151 = node150_l;
      node152 = node150_r;
      node153_r = node145_r & pixel[595];
      node153_l = node145_r & ~pixel[595];
      node154_r = node153_l & pixel[289];
      node154_l = node153_l & ~pixel[289];
      node155 = node154_l;
      node156 = node154_r;
      node157_r = node153_r & pixel[357];
      node157_l = node153_r & ~pixel[357];
      node158 = node157_l;
      node159 = node157_r;
      node160_r = node144_r & pixel[317];
      node160_l = node144_r & ~pixel[317];
      node161_r = node160_l & pixel[514];
      node161_l = node160_l & ~pixel[514];
      node162_r = node161_l & pixel[185];
      node162_l = node161_l & ~pixel[185];
      node163 = node162_l;
      node164 = node162_r;
      node165_r = node161_r & pixel[411];
      node165_l = node161_r & ~pixel[411];
      node166 = node165_l;
      node167 = node165_r;
      node168_r = node160_r & pixel[495];
      node168_l = node160_r & ~pixel[495];
      node169_r = node168_l & pixel[146];
      node169_l = node168_l & ~pixel[146];
      node170 = node169_l;
      node171 = node169_r;
      node172_r = node168_r & pixel[234];
      node172_l = node168_r & ~pixel[234];
      node173 = node172_l;
      node174 = node172_r;
      node175_r = node111_r & pixel[397];
      node175_l = node111_r & ~pixel[397];
      node176_r = node175_l & pixel[593];
      node176_l = node175_l & ~pixel[593];
      node177_r = node176_l & pixel[430];
      node177_l = node176_l & ~pixel[430];
      node178_r = node177_l & pixel[379];
      node178_l = node177_l & ~pixel[379];
      node179_r = node178_l & pixel[568];
      node179_l = node178_l & ~pixel[568];
      node180 = node179_l;
      node181 = node179_r;
      node182_r = node178_r & pixel[524];
      node182_l = node178_r & ~pixel[524];
      node183 = node182_l;
      node184 = node182_r;
      node185_r = node177_r & pixel[123];
      node185_l = node177_r & ~pixel[123];
      node186_r = node185_l & pixel[298];
      node186_l = node185_l & ~pixel[298];
      node187 = node186_l;
      node188 = node186_r;
      node189_r = node185_r & pixel[438];
      node189_l = node185_r & ~pixel[438];
      node190 = node189_l;
      node191 = node189_r;
      node192_r = node176_r & pixel[570];
      node192_l = node176_r & ~pixel[570];
      node193_r = node192_l & pixel[572];
      node193_l = node192_l & ~pixel[572];
      node194 = node193_l;
      node195_r = node193_r & pixel[189];
      node195_l = node193_r & ~pixel[189];
      node196 = node195_l;
      node197 = node195_r;
      node198 = node192_r;
      node199 = node175_r;
      node200_r = node2_r & pixel[525];
      node200_l = node2_r & ~pixel[525];
      node201_r = node200_l & pixel[290];
      node201_l = node200_l & ~pixel[290];
      node202_r = node201_l & pixel[157];
      node202_l = node201_l & ~pixel[157];
      node203_r = node202_l & pixel[635];
      node203_l = node202_l & ~pixel[635];
      node204_r = node203_l & pixel[516];
      node204_l = node203_l & ~pixel[516];
      node205_r = node204_l & pixel[152];
      node205_l = node204_l & ~pixel[152];
      node206_r = node205_l & pixel[372];
      node206_l = node205_l & ~pixel[372];
      node207 = node206_l;
      node208 = node206_r;
      node209_r = node205_r & pixel[489];
      node209_l = node205_r & ~pixel[489];
      node210 = node209_l;
      node211 = node209_r;
      node212_r = node204_r & pixel[541];
      node212_l = node204_r & ~pixel[541];
      node213_r = node212_l & pixel[546];
      node213_l = node212_l & ~pixel[546];
      node214 = node213_l;
      node215 = node213_r;
      node216_r = node212_r & pixel[528];
      node216_l = node212_r & ~pixel[528];
      node217 = node216_l;
      node218 = node216_r;
      node219_r = node203_r & pixel[181];
      node219_l = node203_r & ~pixel[181];
      node220_r = node219_l & pixel[238];
      node220_l = node219_l & ~pixel[238];
      node221_r = node220_l & pixel[180];
      node221_l = node220_l & ~pixel[180];
      node222 = node221_l;
      node223 = node221_r;
      node224_r = node220_r & pixel[379];
      node224_l = node220_r & ~pixel[379];
      node225 = node224_l;
      node226 = node224_r;
      node227_r = node219_r & pixel[456];
      node227_l = node219_r & ~pixel[456];
      node228_r = node227_l & pixel[322];
      node228_l = node227_l & ~pixel[322];
      node229 = node228_l;
      node230 = node228_r;
      node231_r = node227_r & pixel[467];
      node231_l = node227_r & ~pixel[467];
      node232 = node231_l;
      node233 = node231_r;
      node234_r = node202_r & pixel[554];
      node234_l = node202_r & ~pixel[554];
      node235_r = node234_l & pixel[627];
      node235_l = node234_l & ~pixel[627];
      node236_r = node235_l & pixel[354];
      node236_l = node235_l & ~pixel[354];
      node237 = node236_l;
      node238_r = node236_r & pixel[314];
      node238_l = node236_r & ~pixel[314];
      node239 = node238_l;
      node240 = node238_r;
      node241_r = node235_r & pixel[323];
      node241_l = node235_r & ~pixel[323];
      node242 = node241_l;
      node243 = node241_r;
      node244_r = node234_r & pixel[351];
      node244_l = node234_r & ~pixel[351];
      node245_r = node244_l & pixel[519];
      node245_l = node244_l & ~pixel[519];
      node246 = node245_l;
      node247 = node245_r;
      node248 = node244_r;
      node249_r = node201_r & pixel[150];
      node249_l = node201_r & ~pixel[150];
      node250_r = node249_l & pixel[178];
      node250_l = node249_l & ~pixel[178];
      node251_r = node250_l & pixel[749];
      node251_l = node250_l & ~pixel[749];
      node252_r = node251_l & pixel[192];
      node252_l = node251_l & ~pixel[192];
      node253_r = node252_l & pixel[510];
      node253_l = node252_l & ~pixel[510];
      node254 = node253_l;
      node255 = node253_r;
      node256 = node252_r;
      node257_r = node251_r & pixel[516];
      node257_l = node251_r & ~pixel[516];
      node258 = node257_l;
      node259 = node257_r;
      node260_r = node250_r & pixel[347];
      node260_l = node250_r & ~pixel[347];
      node261_r = node260_l & pixel[461];
      node261_l = node260_l & ~pixel[461];
      node262_r = node261_l & pixel[455];
      node262_l = node261_l & ~pixel[455];
      node263 = node262_l;
      node264 = node262_r;
      node265 = node261_r;
      node266 = node260_r;
      node267_r = node249_r & pixel[400];
      node267_l = node249_r & ~pixel[400];
      node268 = node267_l;
      node269_r = node267_r & pixel[188];
      node269_l = node267_r & ~pixel[188];
      node270 = node269_l;
      node271 = node269_r;
      node272_r = node200_r & pixel[404];
      node272_l = node200_r & ~pixel[404];
      node273_r = node272_l & pixel[319];
      node273_l = node272_l & ~pixel[319];
      node274_r = node273_l & pixel[427];
      node274_l = node273_l & ~pixel[427];
      node275_r = node274_l & pixel[511];
      node275_l = node274_l & ~pixel[511];
      node276_r = node275_l & pixel[601];
      node276_l = node275_l & ~pixel[601];
      node277_r = node276_l & pixel[288];
      node277_l = node276_l & ~pixel[288];
      node278 = node277_l;
      node279 = node277_r;
      node280_r = node276_r & pixel[741];
      node280_l = node276_r & ~pixel[741];
      node281 = node280_l;
      node282 = node280_r;
      node283_r = node275_r & pixel[579];
      node283_l = node275_r & ~pixel[579];
      node284_r = node283_l & pixel[323];
      node284_l = node283_l & ~pixel[323];
      node285 = node284_l;
      node286 = node284_r;
      node287_r = node283_r & pixel[298];
      node287_l = node283_r & ~pixel[298];
      node288 = node287_l;
      node289 = node287_r;
      node290_r = node274_r & pixel[471];
      node290_l = node274_r & ~pixel[471];
      node291_r = node290_l & pixel[157];
      node291_l = node290_l & ~pixel[157];
      node292_r = node291_l & pixel[273];
      node292_l = node291_l & ~pixel[273];
      node293 = node292_l;
      node294 = node292_r;
      node295 = node291_r;
      node296_r = node290_r & pixel[92];
      node296_l = node290_r & ~pixel[92];
      node297_r = node296_l & pixel[210];
      node297_l = node296_l & ~pixel[210];
      node298 = node297_l;
      node299 = node297_r;
      node300_r = node296_r & pixel[409];
      node300_l = node296_r & ~pixel[409];
      node301 = node300_l;
      node302 = node300_r;
      node303_r = node273_r & pixel[209];
      node303_l = node273_r & ~pixel[209];
      node304_r = node303_l & pixel[523];
      node304_l = node303_l & ~pixel[523];
      node305_r = node304_l & pixel[176];
      node305_l = node304_l & ~pixel[176];
      node306 = node305_l;
      node307 = node305_r;
      node308_r = node304_r & pixel[383];
      node308_l = node304_r & ~pixel[383];
      node309_r = node308_l & pixel[513];
      node309_l = node308_l & ~pixel[513];
      node310 = node309_l;
      node311 = node309_r;
      node312_r = node308_r & pixel[256];
      node312_l = node308_r & ~pixel[256];
      node313 = node312_l;
      node314 = node312_r;
      node315_r = node303_r & pixel[357];
      node315_l = node303_r & ~pixel[357];
      node316_r = node315_l & pixel[690];
      node316_l = node315_l & ~pixel[690];
      node317_r = node316_l & pixel[204];
      node317_l = node316_l & ~pixel[204];
      node318 = node317_l;
      node319 = node317_r;
      node320_r = node316_r & pixel[200];
      node320_l = node316_r & ~pixel[200];
      node321 = node320_l;
      node322 = node320_r;
      node323_r = node315_r & pixel[153];
      node323_l = node315_r & ~pixel[153];
      node324_r = node323_l & pixel[496];
      node324_l = node323_l & ~pixel[496];
      node325 = node324_l;
      node326 = node324_r;
      node327_r = node323_r & pixel[313];
      node327_l = node323_r & ~pixel[313];
      node328 = node327_l;
      node329 = node327_r;
      node330_r = node272_r & pixel[315];
      node330_l = node272_r & ~pixel[315];
      node331_r = node330_l & pixel[301];
      node331_l = node330_l & ~pixel[301];
      node332_r = node331_l & pixel[666];
      node332_l = node331_l & ~pixel[666];
      node333_r = node332_l & pixel[488];
      node333_l = node332_l & ~pixel[488];
      node334_r = node333_l & pixel[371];
      node334_l = node333_l & ~pixel[371];
      node335 = node334_l;
      node336 = node334_r;
      node337 = node333_r;
      node338_r = node332_r & pixel[153];
      node338_l = node332_r & ~pixel[153];
      node339 = node338_l;
      node340 = node338_r;
      node341 = node331_r;
      node342_r = node330_r & pixel[491];
      node342_l = node330_r & ~pixel[491];
      node343_r = node342_l & pixel[515];
      node343_l = node342_l & ~pixel[515];
      node344_r = node343_l & pixel[637];
      node344_l = node343_l & ~pixel[637];
      node345_r = node344_l & pixel[608];
      node345_l = node344_l & ~pixel[608];
      node346 = node345_l;
      node347 = node345_r;
      node348 = node344_r;
      node349_r = node343_r & pixel[326];
      node349_l = node343_r & ~pixel[326];
      node350 = node349_l;
      node351_r = node349_r & pixel[662];
      node351_l = node349_r & ~pixel[662];
      node352 = node351_l;
      node353 = node351_r;
      node354_r = node342_r & pixel[208];
      node354_l = node342_r & ~pixel[208];
      node355 = node354_l;
      node356_r = node354_r & pixel[240];
      node356_l = node354_r & ~pixel[240];
      node357 = node356_l;
      node358 = node356_r;
      node359_r = node1_r & pixel[350];
      node359_l = node1_r & ~pixel[350];
      node360_r = node359_l & pixel[211];
      node360_l = node359_l & ~pixel[211];
      node361_r = node360_l & pixel[464];
      node361_l = node360_l & ~pixel[464];
      node362_r = node361_l & pixel[515];
      node362_l = node361_l & ~pixel[515];
      node363_r = node362_l & pixel[601];
      node363_l = node362_l & ~pixel[601];
      node364_r = node363_l & pixel[156];
      node364_l = node363_l & ~pixel[156];
      node365_r = node364_l & pixel[490];
      node365_l = node364_l & ~pixel[490];
      node366_r = node365_l & pixel[584];
      node366_l = node365_l & ~pixel[584];
      node367 = node366_l;
      node368 = node366_r;
      node369_r = node365_r & pixel[430];
      node369_l = node365_r & ~pixel[430];
      node370 = node369_l;
      node371 = node369_r;
      node372_r = node364_r & pixel[485];
      node372_l = node364_r & ~pixel[485];
      node373_r = node372_l & pixel[285];
      node373_l = node372_l & ~pixel[285];
      node374 = node373_l;
      node375 = node373_r;
      node376_r = node372_r & pixel[597];
      node376_l = node372_r & ~pixel[597];
      node377 = node376_l;
      node378 = node376_r;
      node379_r = node363_r & pixel[654];
      node379_l = node363_r & ~pixel[654];
      node380_r = node379_l & pixel[541];
      node380_l = node379_l & ~pixel[541];
      node381_r = node380_l & pixel[544];
      node381_l = node380_l & ~pixel[544];
      node382 = node381_l;
      node383 = node381_r;
      node384_r = node380_r & pixel[659];
      node384_l = node380_r & ~pixel[659];
      node385 = node384_l;
      node386 = node384_r;
      node387_r = node379_r & pixel[203];
      node387_l = node379_r & ~pixel[203];
      node388_r = node387_l & pixel[708];
      node388_l = node387_l & ~pixel[708];
      node389 = node388_l;
      node390 = node388_r;
      node391 = node387_r;
      node392_r = node362_r & pixel[656];
      node392_l = node362_r & ~pixel[656];
      node393_r = node392_l & pixel[597];
      node393_l = node392_l & ~pixel[597];
      node394_r = node393_l & pixel[323];
      node394_l = node393_l & ~pixel[323];
      node395_r = node394_l & pixel[300];
      node395_l = node394_l & ~pixel[300];
      node396 = node395_l;
      node397 = node395_r;
      node398_r = node394_r & pixel[513];
      node398_l = node394_r & ~pixel[513];
      node399 = node398_l;
      node400 = node398_r;
      node401_r = node393_r & pixel[441];
      node401_l = node393_r & ~pixel[441];
      node402_r = node401_l & pixel[602];
      node402_l = node401_l & ~pixel[602];
      node403 = node402_l;
      node404 = node402_r;
      node405_r = node401_r & pixel[550];
      node405_l = node401_r & ~pixel[550];
      node406 = node405_l;
      node407 = node405_r;
      node408_r = node392_r & pixel[635];
      node408_l = node392_r & ~pixel[635];
      node409_r = node408_l & pixel[382];
      node409_l = node408_l & ~pixel[382];
      node410_r = node409_l & pixel[242];
      node410_l = node409_l & ~pixel[242];
      node411 = node410_l;
      node412 = node410_r;
      node413_r = node409_r & pixel[426];
      node413_l = node409_r & ~pixel[426];
      node414 = node413_l;
      node415 = node413_r;
      node416_r = node408_r & pixel[410];
      node416_l = node408_r & ~pixel[410];
      node417 = node416_l;
      node418_r = node416_r & pixel[346];
      node418_l = node416_r & ~pixel[346];
      node419 = node418_l;
      node420 = node418_r;
      node421_r = node361_r & pixel[552];
      node421_l = node361_r & ~pixel[552];
      node422_r = node421_l & pixel[430];
      node422_l = node421_l & ~pixel[430];
      node423_r = node422_l & pixel[267];
      node423_l = node422_l & ~pixel[267];
      node424_r = node423_l & pixel[182];
      node424_l = node423_l & ~pixel[182];
      node425_r = node424_l & pixel[345];
      node425_l = node424_l & ~pixel[345];
      node426 = node425_l;
      node427 = node425_r;
      node428_r = node424_r & pixel[569];
      node428_l = node424_r & ~pixel[569];
      node429 = node428_l;
      node430 = node428_r;
      node431_r = node423_r & pixel[353];
      node431_l = node423_r & ~pixel[353];
      node432_r = node431_l & pixel[287];
      node432_l = node431_l & ~pixel[287];
      node433 = node432_l;
      node434 = node432_r;
      node435_r = node431_r & pixel[262];
      node435_l = node431_r & ~pixel[262];
      node436 = node435_l;
      node437 = node435_r;
      node438_r = node422_r & pixel[99];
      node438_l = node422_r & ~pixel[99];
      node439_r = node438_l & pixel[381];
      node439_l = node438_l & ~pixel[381];
      node440_r = node439_l & pixel[382];
      node440_l = node439_l & ~pixel[382];
      node441 = node440_l;
      node442 = node440_r;
      node443_r = node439_r & pixel[229];
      node443_l = node439_r & ~pixel[229];
      node444 = node443_l;
      node445 = node443_r;
      node446_r = node438_r & pixel[208];
      node446_l = node438_r & ~pixel[208];
      node447_r = node446_l & pixel[292];
      node447_l = node446_l & ~pixel[292];
      node448 = node447_l;
      node449 = node447_r;
      node450_r = node446_r & pixel[243];
      node450_l = node446_r & ~pixel[243];
      node451 = node450_l;
      node452 = node450_r;
      node453_r = node421_r & pixel[543];
      node453_l = node421_r & ~pixel[543];
      node454_r = node453_l & pixel[154];
      node454_l = node453_l & ~pixel[154];
      node455_r = node454_l & pixel[599];
      node455_l = node454_l & ~pixel[599];
      node456_r = node455_l & pixel[238];
      node456_l = node455_l & ~pixel[238];
      node457 = node456_l;
      node458 = node456_r;
      node459_r = node455_r & pixel[630];
      node459_l = node455_r & ~pixel[630];
      node460 = node459_l;
      node461 = node459_r;
      node462_r = node454_r & pixel[442];
      node462_l = node454_r & ~pixel[442];
      node463_r = node462_l & pixel[382];
      node463_l = node462_l & ~pixel[382];
      node464 = node463_l;
      node465 = node463_r;
      node466_r = node462_r & pixel[487];
      node466_l = node462_r & ~pixel[487];
      node467 = node466_l;
      node468 = node466_r;
      node469_r = node453_r & pixel[486];
      node469_l = node453_r & ~pixel[486];
      node470_r = node469_l & pixel[659];
      node470_l = node469_l & ~pixel[659];
      node471_r = node470_l & pixel[599];
      node471_l = node470_l & ~pixel[599];
      node472 = node471_l;
      node473 = node471_r;
      node474_r = node470_r & pixel[271];
      node474_l = node470_r & ~pixel[271];
      node475 = node474_l;
      node476 = node474_r;
      node477_r = node469_r & pixel[578];
      node477_l = node469_r & ~pixel[578];
      node478_r = node477_l & pixel[398];
      node478_l = node477_l & ~pixel[398];
      node479 = node478_l;
      node480 = node478_r;
      node481_r = node477_r & pixel[217];
      node481_l = node477_r & ~pixel[217];
      node482 = node481_l;
      node483 = node481_r;
      node484_r = node360_r & pixel[102];
      node484_l = node360_r & ~pixel[102];
      node485_r = node484_l & pixel[542];
      node485_l = node484_l & ~pixel[542];
      node486_r = node485_l & pixel[161];
      node486_l = node485_l & ~pixel[161];
      node487_r = node486_l & pixel[326];
      node487_l = node486_l & ~pixel[326];
      node488_r = node487_l & pixel[653];
      node488_l = node487_l & ~pixel[653];
      node489_r = node488_l & pixel[217];
      node489_l = node488_l & ~pixel[217];
      node490 = node489_l;
      node491 = node489_r;
      node492_r = node488_r & pixel[709];
      node492_l = node488_r & ~pixel[709];
      node493 = node492_l;
      node494 = node492_r;
      node495_r = node487_r & pixel[237];
      node495_l = node487_r & ~pixel[237];
      node496_r = node495_l & pixel[316];
      node496_l = node495_l & ~pixel[316];
      node497 = node496_l;
      node498 = node496_r;
      node499_r = node495_r & pixel[401];
      node499_l = node495_r & ~pixel[401];
      node500 = node499_l;
      node501 = node499_r;
      node502_r = node486_r & pixel[326];
      node502_l = node486_r & ~pixel[326];
      node503_r = node502_l & pixel[356];
      node503_l = node502_l & ~pixel[356];
      node504_r = node503_l & pixel[217];
      node504_l = node503_l & ~pixel[217];
      node505 = node504_l;
      node506 = node504_r;
      node507_r = node503_r & pixel[131];
      node507_l = node503_r & ~pixel[131];
      node508 = node507_l;
      node509 = node507_r;
      node510_r = node502_r & pixel[623];
      node510_l = node502_r & ~pixel[623];
      node511_r = node510_l & pixel[678];
      node511_l = node510_l & ~pixel[678];
      node512 = node511_l;
      node513 = node511_r;
      node514_r = node510_r & pixel[294];
      node514_l = node510_r & ~pixel[294];
      node515 = node514_l;
      node516 = node514_r;
      node517_r = node485_r & pixel[683];
      node517_l = node485_r & ~pixel[683];
      node518_r = node517_l & pixel[325];
      node518_l = node517_l & ~pixel[325];
      node519_r = node518_l & pixel[215];
      node519_l = node518_l & ~pixel[215];
      node520_r = node519_l & pixel[574];
      node520_l = node519_l & ~pixel[574];
      node521 = node520_l;
      node522 = node520_r;
      node523_r = node519_r & pixel[660];
      node523_l = node519_r & ~pixel[660];
      node524 = node523_l;
      node525 = node523_r;
      node526_r = node518_r & pixel[708];
      node526_l = node518_r & ~pixel[708];
      node527_r = node526_l & pixel[319];
      node527_l = node526_l & ~pixel[319];
      node528 = node527_l;
      node529 = node527_r;
      node530_r = node526_r & pixel[404];
      node530_l = node526_r & ~pixel[404];
      node531 = node530_l;
      node532 = node530_r;
      node533_r = node517_r & pixel[184];
      node533_l = node517_r & ~pixel[184];
      node534_r = node533_l & pixel[376];
      node534_l = node533_l & ~pixel[376];
      node535_r = node534_l & pixel[297];
      node535_l = node534_l & ~pixel[297];
      node536 = node535_l;
      node537 = node535_r;
      node538_r = node534_r & pixel[465];
      node538_l = node534_r & ~pixel[465];
      node539 = node538_l;
      node540 = node538_r;
      node541_r = node533_r & pixel[708];
      node541_l = node533_r & ~pixel[708];
      node542_r = node541_l & pixel[149];
      node542_l = node541_l & ~pixel[149];
      node543 = node542_l;
      node544 = node542_r;
      node545_r = node541_r & pixel[374];
      node545_l = node541_r & ~pixel[374];
      node546 = node545_l;
      node547 = node545_r;
      node548_r = node484_r & pixel[481];
      node548_l = node484_r & ~pixel[481];
      node549_r = node548_l & pixel[467];
      node549_l = node548_l & ~pixel[467];
      node550_r = node549_l & pixel[324];
      node550_l = node549_l & ~pixel[324];
      node551_r = node550_l & pixel[484];
      node551_l = node550_l & ~pixel[484];
      node552_r = node551_l & pixel[515];
      node552_l = node551_l & ~pixel[515];
      node553 = node552_l;
      node554 = node552_r;
      node555 = node551_r;
      node556_r = node550_r & pixel[354];
      node556_l = node550_r & ~pixel[354];
      node557 = node556_l;
      node558 = node556_r;
      node559_r = node549_r & pixel[265];
      node559_l = node549_r & ~pixel[265];
      node560_r = node559_l & pixel[568];
      node560_l = node559_l & ~pixel[568];
      node561 = node560_l;
      node562 = node560_r;
      node563 = node559_r;
      node564 = node548_r;
      node565_r = node359_r & pixel[493];
      node565_l = node359_r & ~pixel[493];
      node566_r = node565_l & pixel[375];
      node566_l = node565_l & ~pixel[375];
      node567_r = node566_l & pixel[207];
      node567_l = node566_l & ~pixel[207];
      node568_r = node567_l & pixel[328];
      node568_l = node567_l & ~pixel[328];
      node569_r = node568_l & pixel[606];
      node569_l = node568_l & ~pixel[606];
      node570_r = node569_l & pixel[345];
      node570_l = node569_l & ~pixel[345];
      node571_r = node570_l & pixel[274];
      node571_l = node570_l & ~pixel[274];
      node572 = node571_l;
      node573 = node571_r;
      node574_r = node570_r & pixel[401];
      node574_l = node570_r & ~pixel[401];
      node575 = node574_l;
      node576 = node574_r;
      node577_r = node569_r & pixel[570];
      node577_l = node569_r & ~pixel[570];
      node578_r = node577_l & pixel[179];
      node578_l = node577_l & ~pixel[179];
      node579 = node578_l;
      node580 = node578_r;
      node581_r = node577_r & pixel[515];
      node581_l = node577_r & ~pixel[515];
      node582 = node581_l;
      node583 = node581_r;
      node584_r = node568_r & pixel[524];
      node584_l = node568_r & ~pixel[524];
      node585_r = node584_l & pixel[210];
      node585_l = node584_l & ~pixel[210];
      node586_r = node585_l & pixel[574];
      node586_l = node585_l & ~pixel[574];
      node587 = node586_l;
      node588 = node586_r;
      node589_r = node585_r & pixel[321];
      node589_l = node585_r & ~pixel[321];
      node590 = node589_l;
      node591 = node589_r;
      node592_r = node584_r & pixel[659];
      node592_l = node584_r & ~pixel[659];
      node593_r = node592_l & pixel[544];
      node593_l = node592_l & ~pixel[544];
      node594 = node593_l;
      node595 = node593_r;
      node596_r = node592_r & pixel[205];
      node596_l = node592_r & ~pixel[205];
      node597 = node596_l;
      node598 = node596_r;
      node599_r = node567_r & pixel[320];
      node599_l = node567_r & ~pixel[320];
      node600_r = node599_l & pixel[318];
      node600_l = node599_l & ~pixel[318];
      node601_r = node600_l & pixel[439];
      node601_l = node600_l & ~pixel[439];
      node602_r = node601_l & pixel[178];
      node602_l = node601_l & ~pixel[178];
      node603 = node602_l;
      node604 = node602_r;
      node605_r = node601_r & pixel[495];
      node605_l = node601_r & ~pixel[495];
      node606 = node605_l;
      node607 = node605_r;
      node608_r = node600_r & pixel[211];
      node608_l = node600_r & ~pixel[211];
      node609_r = node608_l & pixel[578];
      node609_l = node608_l & ~pixel[578];
      node610 = node609_l;
      node611 = node609_r;
      node612_r = node608_r & pixel[528];
      node612_l = node608_r & ~pixel[528];
      node613 = node612_l;
      node614 = node612_r;
      node615_r = node599_r & pixel[543];
      node615_l = node599_r & ~pixel[543];
      node616_r = node615_l & pixel[325];
      node616_l = node615_l & ~pixel[325];
      node617_r = node616_l & pixel[351];
      node617_l = node616_l & ~pixel[351];
      node618 = node617_l;
      node619 = node617_r;
      node620_r = node616_r & pixel[406];
      node620_l = node616_r & ~pixel[406];
      node621 = node620_l;
      node622 = node620_r;
      node623_r = node615_r & pixel[377];
      node623_l = node615_r & ~pixel[377];
      node624_r = node623_l & pixel[231];
      node624_l = node623_l & ~pixel[231];
      node625 = node624_l;
      node626 = node624_r;
      node627_r = node623_r & pixel[118];
      node627_l = node623_r & ~pixel[118];
      node628 = node627_l;
      node629 = node627_r;
      node630_r = node566_r & pixel[517];
      node630_l = node566_r & ~pixel[517];
      node631_r = node630_l & pixel[542];
      node631_l = node630_l & ~pixel[542];
      node632_r = node631_l & pixel[492];
      node632_l = node631_l & ~pixel[492];
      node633_r = node632_l & pixel[369];
      node633_l = node632_l & ~pixel[369];
      node634_r = node633_l & pixel[261];
      node634_l = node633_l & ~pixel[261];
      node635 = node634_l;
      node636 = node634_r;
      node637_r = node633_r & pixel[323];
      node637_l = node633_r & ~pixel[323];
      node638 = node637_l;
      node639 = node637_r;
      node640_r = node632_r & pixel[236];
      node640_l = node632_r & ~pixel[236];
      node641_r = node640_l & pixel[268];
      node641_l = node640_l & ~pixel[268];
      node642 = node641_l;
      node643 = node641_r;
      node644_r = node640_r & pixel[179];
      node644_l = node640_r & ~pixel[179];
      node645 = node644_l;
      node646 = node644_r;
      node647_r = node631_r & pixel[215];
      node647_l = node631_r & ~pixel[215];
      node648_r = node647_l & pixel[243];
      node648_l = node647_l & ~pixel[243];
      node649_r = node648_l & pixel[178];
      node649_l = node648_l & ~pixel[178];
      node650 = node649_l;
      node651 = node649_r;
      node652_r = node648_r & pixel[407];
      node652_l = node648_r & ~pixel[407];
      node653 = node652_l;
      node654 = node652_r;
      node655_r = node647_r & pixel[519];
      node655_l = node647_r & ~pixel[519];
      node656_r = node655_l & pixel[574];
      node656_l = node655_l & ~pixel[574];
      node657 = node656_l;
      node658 = node656_r;
      node659_r = node655_r & pixel[105];
      node659_l = node655_r & ~pixel[105];
      node660 = node659_l;
      node661 = node659_r;
      node662_r = node630_r & pixel[606];
      node662_l = node630_r & ~pixel[606];
      node663_r = node662_l & pixel[413];
      node663_l = node662_l & ~pixel[413];
      node664_r = node663_l & pixel[354];
      node664_l = node663_l & ~pixel[354];
      node665_r = node664_l & pixel[243];
      node665_l = node664_l & ~pixel[243];
      node666 = node665_l;
      node667 = node665_r;
      node668_r = node664_r & pixel[155];
      node668_l = node664_r & ~pixel[155];
      node669 = node668_l;
      node670 = node668_r;
      node671_r = node663_r & pixel[524];
      node671_l = node663_r & ~pixel[524];
      node672_r = node671_l & pixel[287];
      node672_l = node671_l & ~pixel[287];
      node673 = node672_l;
      node674 = node672_r;
      node675_r = node671_r & pixel[628];
      node675_l = node671_r & ~pixel[628];
      node676 = node675_l;
      node677 = node675_r;
      node678_r = node662_r & pixel[575];
      node678_l = node662_r & ~pixel[575];
      node679_r = node678_l & pixel[633];
      node679_l = node678_l & ~pixel[633];
      node680 = node679_l;
      node681_r = node679_r & pixel[569];
      node681_l = node679_r & ~pixel[569];
      node682 = node681_l;
      node683 = node681_r;
      node684_r = node678_r & pixel[242];
      node684_l = node678_r & ~pixel[242];
      node685_r = node684_l & pixel[458];
      node685_l = node684_l & ~pixel[458];
      node686 = node685_l;
      node687 = node685_r;
      node688_r = node684_r & pixel[106];
      node688_l = node684_r & ~pixel[106];
      node689 = node688_l;
      node690 = node688_r;
      node691_r = node565_r & pixel[655];
      node691_l = node565_r & ~pixel[655];
      node692_r = node691_l & pixel[400];
      node692_l = node691_l & ~pixel[400];
      node693_r = node692_l & pixel[660];
      node693_l = node692_l & ~pixel[660];
      node694_r = node693_l & pixel[204];
      node694_l = node693_l & ~pixel[204];
      node695_r = node694_l & pixel[542];
      node695_l = node694_l & ~pixel[542];
      node696_r = node695_l & pixel[516];
      node696_l = node695_l & ~pixel[516];
      node697 = node696_l;
      node698 = node696_r;
      node699_r = node695_r & pixel[574];
      node699_l = node695_r & ~pixel[574];
      node700 = node699_l;
      node701 = node699_r;
      node702_r = node694_r & pixel[524];
      node702_l = node694_r & ~pixel[524];
      node703_r = node702_l & pixel[689];
      node703_l = node702_l & ~pixel[689];
      node704 = node703_l;
      node705 = node703_r;
      node706_r = node702_r & pixel[605];
      node706_l = node702_r & ~pixel[605];
      node707 = node706_l;
      node708 = node706_r;
      node709_r = node693_r & pixel[547];
      node709_l = node693_r & ~pixel[547];
      node710_r = node709_l & pixel[488];
      node710_l = node709_l & ~pixel[488];
      node711_r = node710_l & pixel[158];
      node711_l = node710_l & ~pixel[158];
      node712 = node711_l;
      node713 = node711_r;
      node714_r = node710_r & pixel[712];
      node714_l = node710_r & ~pixel[712];
      node715 = node714_l;
      node716 = node714_r;
      node717_r = node709_r & pixel[203];
      node717_l = node709_r & ~pixel[203];
      node718_r = node717_l & pixel[317];
      node718_l = node717_l & ~pixel[317];
      node719 = node718_l;
      node720 = node718_r;
      node721_r = node717_r & pixel[715];
      node721_l = node717_r & ~pixel[715];
      node722 = node721_l;
      node723 = node721_r;
      node724_r = node692_r & pixel[573];
      node724_l = node692_r & ~pixel[573];
      node725_r = node724_l & pixel[742];
      node725_l = node724_l & ~pixel[742];
      node726_r = node725_l & pixel[525];
      node726_l = node725_l & ~pixel[525];
      node727_r = node726_l & pixel[215];
      node727_l = node726_l & ~pixel[215];
      node728 = node727_l;
      node729 = node727_r;
      node730_r = node726_r & pixel[454];
      node730_l = node726_r & ~pixel[454];
      node731 = node730_l;
      node732 = node730_r;
      node733_r = node725_r & pixel[381];
      node733_l = node725_r & ~pixel[381];
      node734_r = node733_l & pixel[352];
      node734_l = node733_l & ~pixel[352];
      node735 = node734_l;
      node736 = node734_r;
      node737_r = node733_r & pixel[357];
      node737_l = node733_r & ~pixel[357];
      node738 = node737_l;
      node739 = node737_r;
      node740_r = node724_r & pixel[544];
      node740_l = node724_r & ~pixel[544];
      node741_r = node740_l & pixel[236];
      node741_l = node740_l & ~pixel[236];
      node742_r = node741_l & pixel[566];
      node742_l = node741_l & ~pixel[566];
      node743 = node742_l;
      node744 = node742_r;
      node745_r = node741_r & pixel[626];
      node745_l = node741_r & ~pixel[626];
      node746 = node745_l;
      node747 = node745_r;
      node748_r = node740_r & pixel[268];
      node748_l = node740_r & ~pixel[268];
      node749_r = node748_l & pixel[245];
      node749_l = node748_l & ~pixel[245];
      node750 = node749_l;
      node751 = node749_r;
      node752_r = node748_r & pixel[261];
      node752_l = node748_r & ~pixel[261];
      node753 = node752_l;
      node754 = node752_r;
      node755_r = node691_r & pixel[486];
      node755_l = node691_r & ~pixel[486];
      node756_r = node755_l & pixel[514];
      node756_l = node755_l & ~pixel[514];
      node757_r = node756_l & pixel[264];
      node757_l = node756_l & ~pixel[264];
      node758_r = node757_l & pixel[544];
      node758_l = node757_l & ~pixel[544];
      node759_r = node758_l & pixel[181];
      node759_l = node758_l & ~pixel[181];
      node760 = node759_l;
      node761 = node759_r;
      node762_r = node758_r & pixel[461];
      node762_l = node758_r & ~pixel[461];
      node763 = node762_l;
      node764 = node762_r;
      node765_r = node757_r & pixel[159];
      node765_l = node757_r & ~pixel[159];
      node766_r = node765_l & pixel[327];
      node766_l = node765_l & ~pixel[327];
      node767 = node766_l;
      node768 = node766_r;
      node769_r = node765_r & pixel[318];
      node769_l = node765_r & ~pixel[318];
      node770 = node769_l;
      node771 = node769_r;
      node772_r = node756_r & pixel[403];
      node772_l = node756_r & ~pixel[403];
      node773_r = node772_l & pixel[290];
      node773_l = node772_l & ~pixel[290];
      node774_r = node773_l & pixel[472];
      node774_l = node773_l & ~pixel[472];
      node775 = node774_l;
      node776 = node774_r;
      node777_r = node773_r & pixel[580];
      node777_l = node773_r & ~pixel[580];
      node778 = node777_l;
      node779 = node777_r;
      node780_r = node772_r & pixel[176];
      node780_l = node772_r & ~pixel[176];
      node781_r = node780_l & pixel[685];
      node781_l = node780_l & ~pixel[685];
      node782 = node781_l;
      node783 = node781_r;
      node784_r = node780_r & pixel[317];
      node784_l = node780_r & ~pixel[317];
      node785 = node784_l;
      node786 = node784_r;
      node787_r = node755_r & pixel[430];
      node787_l = node755_r & ~pixel[430];
      node788_r = node787_l & pixel[657];
      node788_l = node787_l & ~pixel[657];
      node789_r = node788_l & pixel[159];
      node789_l = node788_l & ~pixel[159];
      node790_r = node789_l & pixel[522];
      node790_l = node789_l & ~pixel[522];
      node791 = node790_l;
      node792 = node790_r;
      node793_r = node789_r & pixel[183];
      node793_l = node789_r & ~pixel[183];
      node794 = node793_l;
      node795 = node793_r;
      node796_r = node788_r & pixel[484];
      node796_l = node788_r & ~pixel[484];
      node797_r = node796_l & pixel[442];
      node797_l = node796_l & ~pixel[442];
      node798 = node797_l;
      node799 = node797_r;
      node800_r = node796_r & pixel[524];
      node800_l = node796_r & ~pixel[524];
      node801 = node800_l;
      node802 = node800_r;
      node803_r = node787_r & pixel[513];
      node803_l = node787_r & ~pixel[513];
      node804_r = node803_l & pixel[372];
      node804_l = node803_l & ~pixel[372];
      node805_r = node804_l & pixel[651];
      node805_l = node804_l & ~pixel[651];
      node806 = node805_l;
      node807 = node805_r;
      node808_r = node804_r & pixel[316];
      node808_l = node804_r & ~pixel[316];
      node809 = node808_l;
      node810 = node808_r;
      node811_r = node803_r & pixel[181];
      node811_l = node803_r & ~pixel[181];
      node812_r = node811_l & pixel[159];
      node812_l = node811_l & ~pixel[159];
      node813 = node812_l;
      node814 = node812_r;
      node815_r = node811_r & pixel[290];
      node815_l = node811_r & ~pixel[290];
      node816 = node815_l;
      node817 = node815_r;
      node818_r = node0_r & pixel[460];
      node818_l = node0_r & ~pixel[460];
      node819_r = node818_l & pixel[329];
      node819_l = node818_l & ~pixel[329];
      node820_r = node819_l & pixel[387];
      node820_l = node819_l & ~pixel[387];
      node821_r = node820_l & pixel[155];
      node821_l = node820_l & ~pixel[155];
      node822_r = node821_l & pixel[327];
      node822_l = node821_l & ~pixel[327];
      node823_r = node822_l & pixel[102];
      node823_l = node822_l & ~pixel[102];
      node824_r = node823_l & pixel[190];
      node824_l = node823_l & ~pixel[190];
      node825_r = node824_l & pixel[158];
      node825_l = node824_l & ~pixel[158];
      node826_r = node825_l & pixel[176];
      node826_l = node825_l & ~pixel[176];
      node827 = node826_l;
      node828 = node826_r;
      node829_r = node825_r & pixel[624];
      node829_l = node825_r & ~pixel[624];
      node830 = node829_l;
      node831 = node829_r;
      node832_r = node824_r & pixel[322];
      node832_l = node824_r & ~pixel[322];
      node833_r = node832_l & pixel[487];
      node833_l = node832_l & ~pixel[487];
      node834 = node833_l;
      node835 = node833_r;
      node836_r = node832_r & pixel[80];
      node836_l = node832_r & ~pixel[80];
      node837 = node836_l;
      node838 = node836_r;
      node839_r = node823_r & pixel[430];
      node839_l = node823_r & ~pixel[430];
      node840_r = node839_l & pixel[295];
      node840_l = node839_l & ~pixel[295];
      node841_r = node840_l & pixel[464];
      node841_l = node840_l & ~pixel[464];
      node842 = node841_l;
      node843 = node841_r;
      node844_r = node840_r & pixel[497];
      node844_l = node840_r & ~pixel[497];
      node845 = node844_l;
      node846 = node844_r;
      node847_r = node839_r & pixel[622];
      node847_l = node839_r & ~pixel[622];
      node848_r = node847_l & pixel[495];
      node848_l = node847_l & ~pixel[495];
      node849 = node848_l;
      node850 = node848_r;
      node851 = node847_r;
      node852_r = node822_r & pixel[248];
      node852_l = node822_r & ~pixel[248];
      node853_r = node852_l & pixel[485];
      node853_l = node852_l & ~pixel[485];
      node854_r = node853_l & pixel[576];
      node854_l = node853_l & ~pixel[576];
      node855_r = node854_l & pixel[465];
      node855_l = node854_l & ~pixel[465];
      node856 = node855_l;
      node857 = node855_r;
      node858_r = node854_r & pixel[300];
      node858_l = node854_r & ~pixel[300];
      node859 = node858_l;
      node860 = node858_r;
      node861_r = node853_r & pixel[570];
      node861_l = node853_r & ~pixel[570];
      node862_r = node861_l & pixel[156];
      node862_l = node861_l & ~pixel[156];
      node863 = node862_l;
      node864 = node862_r;
      node865_r = node861_r & pixel[441];
      node865_l = node861_r & ~pixel[441];
      node866 = node865_l;
      node867 = node865_r;
      node868_r = node852_r & pixel[610];
      node868_l = node852_r & ~pixel[610];
      node869_r = node868_l & pixel[412];
      node869_l = node868_l & ~pixel[412];
      node870_r = node869_l & pixel[276];
      node870_l = node869_l & ~pixel[276];
      node871 = node870_l;
      node872 = node870_r;
      node873 = node869_r;
      node874 = node868_r;
      node875_r = node821_r & pixel[349];
      node875_l = node821_r & ~pixel[349];
      node876_r = node875_l & pixel[292];
      node876_l = node875_l & ~pixel[292];
      node877_r = node876_l & pixel[518];
      node877_l = node876_l & ~pixel[518];
      node878_r = node877_l & pixel[427];
      node878_l = node877_l & ~pixel[427];
      node879_r = node878_l & pixel[162];
      node879_l = node878_l & ~pixel[162];
      node880 = node879_l;
      node881 = node879_r;
      node882_r = node878_r & pixel[431];
      node882_l = node878_r & ~pixel[431];
      node883 = node882_l;
      node884 = node882_r;
      node885_r = node877_r & pixel[410];
      node885_l = node877_r & ~pixel[410];
      node886_r = node885_l & pixel[289];
      node886_l = node885_l & ~pixel[289];
      node887 = node886_l;
      node888 = node886_r;
      node889_r = node885_r & pixel[345];
      node889_l = node885_r & ~pixel[345];
      node890 = node889_l;
      node891 = node889_r;
      node892_r = node876_r & pixel[214];
      node892_l = node876_r & ~pixel[214];
      node893_r = node892_l & pixel[491];
      node893_l = node892_l & ~pixel[491];
      node894_r = node893_l & pixel[544];
      node894_l = node893_l & ~pixel[544];
      node895 = node894_l;
      node896 = node894_r;
      node897_r = node893_r & pixel[128];
      node897_l = node893_r & ~pixel[128];
      node898 = node897_l;
      node899 = node897_r;
      node900_r = node892_r & pixel[160];
      node900_l = node892_r & ~pixel[160];
      node901_r = node900_l & pixel[347];
      node901_l = node900_l & ~pixel[347];
      node902 = node901_l;
      node903 = node901_r;
      node904_r = node900_r & pixel[401];
      node904_l = node900_r & ~pixel[401];
      node905 = node904_l;
      node906 = node904_r;
      node907_r = node875_r & pixel[263];
      node907_l = node875_r & ~pixel[263];
      node908_r = node907_l & pixel[270];
      node908_l = node907_l & ~pixel[270];
      node909_r = node908_l & pixel[190];
      node909_l = node908_l & ~pixel[190];
      node910_r = node909_l & pixel[240];
      node910_l = node909_l & ~pixel[240];
      node911 = node910_l;
      node912 = node910_r;
      node913_r = node909_r & pixel[357];
      node913_l = node909_r & ~pixel[357];
      node914 = node913_l;
      node915 = node913_r;
      node916_r = node908_r & pixel[152];
      node916_l = node908_r & ~pixel[152];
      node917_r = node916_l & pixel[383];
      node917_l = node916_l & ~pixel[383];
      node918 = node917_l;
      node919 = node917_r;
      node920_r = node916_r & pixel[610];
      node920_l = node916_r & ~pixel[610];
      node921 = node920_l;
      node922 = node920_r;
      node923_r = node907_r & pixel[269];
      node923_l = node907_r & ~pixel[269];
      node924_r = node923_l & pixel[458];
      node924_l = node923_l & ~pixel[458];
      node925_r = node924_l & pixel[569];
      node925_l = node924_l & ~pixel[569];
      node926 = node925_l;
      node927 = node925_r;
      node928_r = node924_r & pixel[271];
      node928_l = node924_r & ~pixel[271];
      node929 = node928_l;
      node930 = node928_r;
      node931_r = node923_r & pixel[428];
      node931_l = node923_r & ~pixel[428];
      node932_r = node931_l & pixel[458];
      node932_l = node931_l & ~pixel[458];
      node933 = node932_l;
      node934 = node932_r;
      node935_r = node931_r & pixel[180];
      node935_l = node931_r & ~pixel[180];
      node936 = node935_l;
      node937 = node935_r;
      node938_r = node820_r & pixel[303];
      node938_l = node820_r & ~pixel[303];
      node939_r = node938_l & pixel[547];
      node939_l = node938_l & ~pixel[547];
      node940_r = node939_l & pixel[173];
      node940_l = node939_l & ~pixel[173];
      node941_r = node940_l & pixel[565];
      node941_l = node940_l & ~pixel[565];
      node942_r = node941_l & pixel[377];
      node942_l = node941_l & ~pixel[377];
      node943_r = node942_l & pixel[183];
      node943_l = node942_l & ~pixel[183];
      node944 = node943_l;
      node945 = node943_r;
      node946_r = node942_r & pixel[573];
      node946_l = node942_r & ~pixel[573];
      node947 = node946_l;
      node948 = node946_r;
      node949_r = node941_r & pixel[470];
      node949_l = node941_r & ~pixel[470];
      node950 = node949_l;
      node951_r = node949_r & pixel[296];
      node951_l = node949_r & ~pixel[296];
      node952 = node951_l;
      node953 = node951_r;
      node954 = node940_r;
      node955_r = node939_r & pixel[576];
      node955_l = node939_r & ~pixel[576];
      node956_r = node955_l & pixel[371];
      node956_l = node955_l & ~pixel[371];
      node957_r = node956_l & pixel[215];
      node957_l = node956_l & ~pixel[215];
      node958 = node957_l;
      node959 = node957_r;
      node960_r = node956_r & pixel[211];
      node960_l = node956_r & ~pixel[211];
      node961 = node960_l;
      node962_r = node960_r & pixel[264];
      node962_l = node960_r & ~pixel[264];
      node963 = node962_l;
      node964 = node962_r;
      node965_r = node955_r & pixel[301];
      node965_l = node955_r & ~pixel[301];
      node966_r = node965_l & pixel[441];
      node966_l = node965_l & ~pixel[441];
      node967_r = node966_l & pixel[470];
      node967_l = node966_l & ~pixel[470];
      node968 = node967_l;
      node969 = node967_r;
      node970 = node966_r;
      node971 = node965_r;
      node972_r = node938_r & pixel[65];
      node972_l = node938_r & ~pixel[65];
      node973_r = node972_l & pixel[120];
      node973_l = node972_l & ~pixel[120];
      node974_r = node973_l & pixel[438];
      node974_l = node973_l & ~pixel[438];
      node975_r = node974_l & pixel[131];
      node975_l = node974_l & ~pixel[131];
      node976 = node975_l;
      node977_r = node975_r & pixel[610];
      node977_l = node975_r & ~pixel[610];
      node978 = node977_l;
      node979 = node977_r;
      node980_r = node974_r & pixel[685];
      node980_l = node974_r & ~pixel[685];
      node981_r = node980_l & pixel[609];
      node981_l = node980_l & ~pixel[609];
      node982 = node981_l;
      node983 = node981_r;
      node984 = node980_r;
      node985_r = node973_r & pixel[152];
      node985_l = node973_r & ~pixel[152];
      node986 = node985_l;
      node987 = node985_r;
      node988 = node972_r;
      node989_r = node819_r & pixel[352];
      node989_l = node819_r & ~pixel[352];
      node990_r = node989_l & pixel[658];
      node990_l = node989_l & ~pixel[658];
      node991_r = node990_l & pixel[238];
      node991_l = node990_l & ~pixel[238];
      node992_r = node991_l & pixel[344];
      node992_l = node991_l & ~pixel[344];
      node993_r = node992_l & pixel[596];
      node993_l = node992_l & ~pixel[596];
      node994_r = node993_l & pixel[243];
      node994_l = node993_l & ~pixel[243];
      node995_r = node994_l & pixel[296];
      node995_l = node994_l & ~pixel[296];
      node996 = node995_l;
      node997 = node995_r;
      node998_r = node994_r & pixel[538];
      node998_l = node994_r & ~pixel[538];
      node999 = node998_l;
      node1000 = node998_r;
      node1001_r = node993_r & pixel[410];
      node1001_l = node993_r & ~pixel[410];
      node1002_r = node1001_l & pixel[242];
      node1002_l = node1001_l & ~pixel[242];
      node1003 = node1002_l;
      node1004 = node1002_r;
      node1005_r = node1001_r & pixel[241];
      node1005_l = node1001_r & ~pixel[241];
      node1006 = node1005_l;
      node1007 = node1005_r;
      node1008_r = node992_r & pixel[492];
      node1008_l = node992_r & ~pixel[492];
      node1009_r = node1008_l & pixel[689];
      node1009_l = node1008_l & ~pixel[689];
      node1010_r = node1009_l & pixel[216];
      node1010_l = node1009_l & ~pixel[216];
      node1011 = node1010_l;
      node1012 = node1010_r;
      node1013_r = node1009_r & pixel[566];
      node1013_l = node1009_r & ~pixel[566];
      node1014 = node1013_l;
      node1015 = node1013_r;
      node1016_r = node1008_r & pixel[212];
      node1016_l = node1008_r & ~pixel[212];
      node1017_r = node1016_l & pixel[273];
      node1017_l = node1016_l & ~pixel[273];
      node1018 = node1017_l;
      node1019 = node1017_r;
      node1020_r = node1016_r & pixel[435];
      node1020_l = node1016_r & ~pixel[435];
      node1021 = node1020_l;
      node1022 = node1020_r;
      node1023_r = node991_r & pixel[73];
      node1023_l = node991_r & ~pixel[73];
      node1024_r = node1023_l & pixel[664];
      node1024_l = node1023_l & ~pixel[664];
      node1025_r = node1024_l & pixel[409];
      node1025_l = node1024_l & ~pixel[409];
      node1026_r = node1025_l & pixel[311];
      node1026_l = node1025_l & ~pixel[311];
      node1027 = node1026_l;
      node1028 = node1026_r;
      node1029_r = node1025_r & pixel[374];
      node1029_l = node1025_r & ~pixel[374];
      node1030 = node1029_l;
      node1031 = node1029_r;
      node1032_r = node1024_r & pixel[376];
      node1032_l = node1024_r & ~pixel[376];
      node1033_r = node1032_l & pixel[410];
      node1033_l = node1032_l & ~pixel[410];
      node1034 = node1033_l;
      node1035 = node1033_r;
      node1036 = node1032_r;
      node1037 = node1023_r;
      node1038_r = node990_r & pixel[378];
      node1038_l = node990_r & ~pixel[378];
      node1039_r = node1038_l & pixel[462];
      node1039_l = node1038_l & ~pixel[462];
      node1040_r = node1039_l & pixel[283];
      node1040_l = node1039_l & ~pixel[283];
      node1041_r = node1040_l & pixel[177];
      node1041_l = node1040_l & ~pixel[177];
      node1042_r = node1041_l & pixel[381];
      node1042_l = node1041_l & ~pixel[381];
      node1043 = node1042_l;
      node1044 = node1042_r;
      node1045_r = node1041_r & pixel[492];
      node1045_l = node1041_r & ~pixel[492];
      node1046 = node1045_l;
      node1047 = node1045_r;
      node1048 = node1040_r;
      node1049_r = node1039_r & pixel[238];
      node1049_l = node1039_r & ~pixel[238];
      node1050_r = node1049_l & pixel[684];
      node1050_l = node1049_l & ~pixel[684];
      node1051 = node1050_l;
      node1052_r = node1050_r & pixel[184];
      node1052_l = node1050_r & ~pixel[184];
      node1053 = node1052_l;
      node1054 = node1052_r;
      node1055_r = node1049_r & pixel[208];
      node1055_l = node1049_r & ~pixel[208];
      node1056 = node1055_l;
      node1057 = node1055_r;
      node1058_r = node1038_r & pixel[463];
      node1058_l = node1038_r & ~pixel[463];
      node1059_r = node1058_l & pixel[654];
      node1059_l = node1058_l & ~pixel[654];
      node1060_r = node1059_l & pixel[656];
      node1060_l = node1059_l & ~pixel[656];
      node1061 = node1060_l;
      node1062 = node1060_r;
      node1063_r = node1059_r & pixel[243];
      node1063_l = node1059_r & ~pixel[243];
      node1064_r = node1063_l & pixel[432];
      node1064_l = node1063_l & ~pixel[432];
      node1065 = node1064_l;
      node1066 = node1064_r;
      node1067 = node1063_r;
      node1068_r = node1058_r & pixel[573];
      node1068_l = node1058_r & ~pixel[573];
      node1069 = node1068_l;
      node1070_r = node1068_r & pixel[466];
      node1070_l = node1068_r & ~pixel[466];
      node1071 = node1070_l;
      node1072_r = node1070_r & pixel[472];
      node1072_l = node1070_r & ~pixel[472];
      node1073 = node1072_l;
      node1074 = node1072_r;
      node1075_r = node989_r & pixel[432];
      node1075_l = node989_r & ~pixel[432];
      node1076_r = node1075_l & pixel[290];
      node1076_l = node1075_l & ~pixel[290];
      node1077_r = node1076_l & pixel[626];
      node1077_l = node1076_l & ~pixel[626];
      node1078_r = node1077_l & pixel[410];
      node1078_l = node1077_l & ~pixel[410];
      node1079_r = node1078_l & pixel[625];
      node1079_l = node1078_l & ~pixel[625];
      node1080_r = node1079_l & pixel[595];
      node1080_l = node1079_l & ~pixel[595];
      node1081 = node1080_l;
      node1082 = node1080_r;
      node1083 = node1079_r;
      node1084_r = node1078_r & pixel[400];
      node1084_l = node1078_r & ~pixel[400];
      node1085_r = node1084_l & pixel[385];
      node1085_l = node1084_l & ~pixel[385];
      node1086 = node1085_l;
      node1087 = node1085_r;
      node1088_r = node1084_r & pixel[267];
      node1088_l = node1084_r & ~pixel[267];
      node1089 = node1088_l;
      node1090 = node1088_r;
      node1091_r = node1077_r & pixel[457];
      node1091_l = node1077_r & ~pixel[457];
      node1092_r = node1091_l & pixel[609];
      node1092_l = node1091_l & ~pixel[609];
      node1093_r = node1092_l & pixel[488];
      node1093_l = node1092_l & ~pixel[488];
      node1094 = node1093_l;
      node1095 = node1093_r;
      node1096_r = node1092_r & pixel[266];
      node1096_l = node1092_r & ~pixel[266];
      node1097 = node1096_l;
      node1098 = node1096_r;
      node1099_r = node1091_r & pixel[498];
      node1099_l = node1091_r & ~pixel[498];
      node1100_r = node1099_l & pixel[357];
      node1100_l = node1099_l & ~pixel[357];
      node1101 = node1100_l;
      node1102 = node1100_r;
      node1103 = node1099_r;
      node1104_r = node1076_r & pixel[436];
      node1104_l = node1076_r & ~pixel[436];
      node1105_r = node1104_l & pixel[264];
      node1105_l = node1104_l & ~pixel[264];
      node1106_r = node1105_l & pixel[359];
      node1106_l = node1105_l & ~pixel[359];
      node1107_r = node1106_l & pixel[575];
      node1107_l = node1106_l & ~pixel[575];
      node1108 = node1107_l;
      node1109 = node1107_r;
      node1110_r = node1106_r & pixel[580];
      node1110_l = node1106_r & ~pixel[580];
      node1111 = node1110_l;
      node1112 = node1110_r;
      node1113_r = node1105_r & pixel[270];
      node1113_l = node1105_r & ~pixel[270];
      node1114_r = node1113_l & pixel[244];
      node1114_l = node1113_l & ~pixel[244];
      node1115 = node1114_l;
      node1116 = node1114_r;
      node1117_r = node1113_r & pixel[454];
      node1117_l = node1113_r & ~pixel[454];
      node1118 = node1117_l;
      node1119 = node1117_r;
      node1120_r = node1104_r & pixel[265];
      node1120_l = node1104_r & ~pixel[265];
      node1121_r = node1120_l & pixel[187];
      node1121_l = node1120_l & ~pixel[187];
      node1122_r = node1121_l & pixel[287];
      node1122_l = node1121_l & ~pixel[287];
      node1123 = node1122_l;
      node1124 = node1122_r;
      node1125_r = node1121_r & pixel[121];
      node1125_l = node1121_r & ~pixel[121];
      node1126 = node1125_l;
      node1127 = node1125_r;
      node1128_r = node1120_r & pixel[240];
      node1128_l = node1120_r & ~pixel[240];
      node1129_r = node1128_l & pixel[216];
      node1129_l = node1128_l & ~pixel[216];
      node1130 = node1129_l;
      node1131 = node1129_r;
      node1132_r = node1128_r & pixel[404];
      node1132_l = node1128_r & ~pixel[404];
      node1133 = node1132_l;
      node1134 = node1132_r;
      node1135_r = node1075_r & pixel[536];
      node1135_l = node1075_r & ~pixel[536];
      node1136_r = node1135_l & pixel[543];
      node1136_l = node1135_l & ~pixel[543];
      node1137_r = node1136_l & pixel[290];
      node1137_l = node1136_l & ~pixel[290];
      node1138_r = node1137_l & pixel[494];
      node1138_l = node1137_l & ~pixel[494];
      node1139_r = node1138_l & pixel[661];
      node1139_l = node1138_l & ~pixel[661];
      node1140 = node1139_l;
      node1141 = node1139_r;
      node1142_r = node1138_r & pixel[382];
      node1142_l = node1138_r & ~pixel[382];
      node1143 = node1142_l;
      node1144 = node1142_r;
      node1145_r = node1137_r & pixel[379];
      node1145_l = node1137_r & ~pixel[379];
      node1146 = node1145_l;
      node1147_r = node1145_r & pixel[415];
      node1147_l = node1145_r & ~pixel[415];
      node1148 = node1147_l;
      node1149 = node1147_r;
      node1150_r = node1136_r & pixel[213];
      node1150_l = node1136_r & ~pixel[213];
      node1151_r = node1150_l & pixel[371];
      node1151_l = node1150_l & ~pixel[371];
      node1152_r = node1151_l & pixel[332];
      node1152_l = node1151_l & ~pixel[332];
      node1153 = node1152_l;
      node1154 = node1152_r;
      node1155 = node1151_r;
      node1156_r = node1150_r & pixel[319];
      node1156_l = node1150_r & ~pixel[319];
      node1157_r = node1156_l & pixel[483];
      node1157_l = node1156_l & ~pixel[483];
      node1158 = node1157_l;
      node1159 = node1157_r;
      node1160_r = node1156_r & pixel[205];
      node1160_l = node1156_r & ~pixel[205];
      node1161 = node1160_l;
      node1162 = node1160_r;
      node1163_r = node1135_r & pixel[326];
      node1163_l = node1135_r & ~pixel[326];
      node1164_r = node1163_l & pixel[692];
      node1164_l = node1163_l & ~pixel[692];
      node1165 = node1164_l;
      node1166 = node1164_r;
      node1167_r = node1163_r & pixel[487];
      node1167_l = node1163_r & ~pixel[487];
      node1168_r = node1167_l & pixel[471];
      node1168_l = node1167_l & ~pixel[471];
      node1169_r = node1168_l & pixel[179];
      node1169_l = node1168_l & ~pixel[179];
      node1170 = node1169_l;
      node1171 = node1169_r;
      node1172 = node1168_r;
      node1173 = node1167_r;
      node1174_r = node818_r & pixel[102];
      node1174_l = node818_r & ~pixel[102];
      node1175_r = node1174_l & pixel[348];
      node1175_l = node1174_l & ~pixel[348];
      node1176_r = node1175_l & pixel[374];
      node1176_l = node1175_l & ~pixel[374];
      node1177_r = node1176_l & pixel[316];
      node1177_l = node1176_l & ~pixel[316];
      node1178_r = node1177_l & pixel[127];
      node1178_l = node1177_l & ~pixel[127];
      node1179_r = node1178_l & pixel[208];
      node1179_l = node1178_l & ~pixel[208];
      node1180_r = node1179_l & pixel[465];
      node1180_l = node1179_l & ~pixel[465];
      node1181_r = node1180_l & pixel[269];
      node1181_l = node1180_l & ~pixel[269];
      node1182 = node1181_l;
      node1183 = node1181_r;
      node1184_r = node1180_r & pixel[271];
      node1184_l = node1180_r & ~pixel[271];
      node1185 = node1184_l;
      node1186 = node1184_r;
      node1187_r = node1179_r & pixel[657];
      node1187_l = node1179_r & ~pixel[657];
      node1188_r = node1187_l & pixel[277];
      node1188_l = node1187_l & ~pixel[277];
      node1189 = node1188_l;
      node1190 = node1188_r;
      node1191_r = node1187_r & pixel[459];
      node1191_l = node1187_r & ~pixel[459];
      node1192 = node1191_l;
      node1193 = node1191_r;
      node1194_r = node1178_r & pixel[97];
      node1194_l = node1178_r & ~pixel[97];
      node1195_r = node1194_l & pixel[396];
      node1195_l = node1194_l & ~pixel[396];
      node1196_r = node1195_l & pixel[516];
      node1196_l = node1195_l & ~pixel[516];
      node1197 = node1196_l;
      node1198 = node1196_r;
      node1199 = node1195_r;
      node1200 = node1194_r;
      node1201_r = node1177_r & pixel[566];
      node1201_l = node1177_r & ~pixel[566];
      node1202_r = node1201_l & pixel[544];
      node1202_l = node1201_l & ~pixel[544];
      node1203_r = node1202_l & pixel[155];
      node1203_l = node1202_l & ~pixel[155];
      node1204_r = node1203_l & pixel[515];
      node1204_l = node1203_l & ~pixel[515];
      node1205 = node1204_l;
      node1206 = node1204_r;
      node1207_r = node1203_r & pixel[385];
      node1207_l = node1203_r & ~pixel[385];
      node1208 = node1207_l;
      node1209 = node1207_r;
      node1210_r = node1202_r & pixel[268];
      node1210_l = node1202_r & ~pixel[268];
      node1211_r = node1210_l & pixel[415];
      node1211_l = node1210_l & ~pixel[415];
      node1212 = node1211_l;
      node1213 = node1211_r;
      node1214_r = node1210_r & pixel[385];
      node1214_l = node1210_r & ~pixel[385];
      node1215 = node1214_l;
      node1216 = node1214_r;
      node1217_r = node1201_r & pixel[545];
      node1217_l = node1201_r & ~pixel[545];
      node1218_r = node1217_l & pixel[486];
      node1218_l = node1217_l & ~pixel[486];
      node1219_r = node1218_l & pixel[381];
      node1219_l = node1218_l & ~pixel[381];
      node1220 = node1219_l;
      node1221 = node1219_r;
      node1222_r = node1218_r & pixel[452];
      node1222_l = node1218_r & ~pixel[452];
      node1223 = node1222_l;
      node1224 = node1222_r;
      node1225_r = node1217_r & pixel[275];
      node1225_l = node1217_r & ~pixel[275];
      node1226_r = node1225_l & pixel[414];
      node1226_l = node1225_l & ~pixel[414];
      node1227 = node1226_l;
      node1228 = node1226_r;
      node1229_r = node1225_r & pixel[604];
      node1229_l = node1225_r & ~pixel[604];
      node1230 = node1229_l;
      node1231 = node1229_r;
      node1232_r = node1176_r & pixel[658];
      node1232_l = node1176_r & ~pixel[658];
      node1233_r = node1232_l & pixel[213];
      node1233_l = node1232_l & ~pixel[213];
      node1234_r = node1233_l & pixel[428];
      node1234_l = node1233_l & ~pixel[428];
      node1235_r = node1234_l & pixel[380];
      node1235_l = node1234_l & ~pixel[380];
      node1236_r = node1235_l & pixel[367];
      node1236_l = node1235_l & ~pixel[367];
      node1237 = node1236_l;
      node1238 = node1236_r;
      node1239_r = node1235_r & pixel[405];
      node1239_l = node1235_r & ~pixel[405];
      node1240 = node1239_l;
      node1241 = node1239_r;
      node1242_r = node1234_r & pixel[187];
      node1242_l = node1234_r & ~pixel[187];
      node1243_r = node1242_l & pixel[574];
      node1243_l = node1242_l & ~pixel[574];
      node1244 = node1243_l;
      node1245 = node1243_r;
      node1246_r = node1242_r & pixel[344];
      node1246_l = node1242_r & ~pixel[344];
      node1247 = node1246_l;
      node1248 = node1246_r;
      node1249_r = node1233_r & pixel[345];
      node1249_l = node1233_r & ~pixel[345];
      node1250_r = node1249_l & pixel[427];
      node1250_l = node1249_l & ~pixel[427];
      node1251_r = node1250_l & pixel[440];
      node1251_l = node1250_l & ~pixel[440];
      node1252 = node1251_l;
      node1253 = node1251_r;
      node1254_r = node1250_r & pixel[340];
      node1254_l = node1250_r & ~pixel[340];
      node1255 = node1254_l;
      node1256 = node1254_r;
      node1257_r = node1249_r & pixel[237];
      node1257_l = node1249_r & ~pixel[237];
      node1258_r = node1257_l & pixel[457];
      node1258_l = node1257_l & ~pixel[457];
      node1259 = node1258_l;
      node1260 = node1258_r;
      node1261_r = node1257_r & pixel[495];
      node1261_l = node1257_r & ~pixel[495];
      node1262 = node1261_l;
      node1263 = node1261_r;
      node1264_r = node1232_r & pixel[595];
      node1264_l = node1232_r & ~pixel[595];
      node1265_r = node1264_l & pixel[156];
      node1265_l = node1264_l & ~pixel[156];
      node1266_r = node1265_l & pixel[293];
      node1266_l = node1265_l & ~pixel[293];
      node1267_r = node1266_l & pixel[493];
      node1267_l = node1266_l & ~pixel[493];
      node1268 = node1267_l;
      node1269 = node1267_r;
      node1270_r = node1266_r & pixel[187];
      node1270_l = node1266_r & ~pixel[187];
      node1271 = node1270_l;
      node1272 = node1270_r;
      node1273_r = node1265_r & pixel[572];
      node1273_l = node1265_r & ~pixel[572];
      node1274_r = node1273_l & pixel[547];
      node1274_l = node1273_l & ~pixel[547];
      node1275 = node1274_l;
      node1276 = node1274_r;
      node1277_r = node1273_r & pixel[383];
      node1277_l = node1273_r & ~pixel[383];
      node1278 = node1277_l;
      node1279 = node1277_r;
      node1280_r = node1264_r & pixel[541];
      node1280_l = node1264_r & ~pixel[541];
      node1281_r = node1280_l & pixel[523];
      node1281_l = node1280_l & ~pixel[523];
      node1282_r = node1281_l & pixel[353];
      node1282_l = node1281_l & ~pixel[353];
      node1283 = node1282_l;
      node1284 = node1282_r;
      node1285_r = node1281_r & pixel[344];
      node1285_l = node1281_r & ~pixel[344];
      node1286 = node1285_l;
      node1287 = node1285_r;
      node1288_r = node1280_r & pixel[408];
      node1288_l = node1280_r & ~pixel[408];
      node1289_r = node1288_l & pixel[270];
      node1289_l = node1288_l & ~pixel[270];
      node1290 = node1289_l;
      node1291 = node1289_r;
      node1292_r = node1288_r & pixel[500];
      node1292_l = node1288_r & ~pixel[500];
      node1293 = node1292_l;
      node1294 = node1292_r;
      node1295_r = node1175_r & pixel[629];
      node1295_l = node1175_r & ~pixel[629];
      node1296_r = node1295_l & pixel[494];
      node1296_l = node1295_l & ~pixel[494];
      node1297_r = node1296_l & pixel[577];
      node1297_l = node1296_l & ~pixel[577];
      node1298_r = node1297_l & pixel[213];
      node1298_l = node1297_l & ~pixel[213];
      node1299_r = node1298_l & pixel[236];
      node1299_l = node1298_l & ~pixel[236];
      node1300_r = node1299_l & pixel[176];
      node1300_l = node1299_l & ~pixel[176];
      node1301 = node1300_l;
      node1302 = node1300_r;
      node1303_r = node1299_r & pixel[162];
      node1303_l = node1299_r & ~pixel[162];
      node1304 = node1303_l;
      node1305 = node1303_r;
      node1306_r = node1298_r & pixel[274];
      node1306_l = node1298_r & ~pixel[274];
      node1307_r = node1306_l & pixel[652];
      node1307_l = node1306_l & ~pixel[652];
      node1308 = node1307_l;
      node1309 = node1307_r;
      node1310_r = node1306_r & pixel[520];
      node1310_l = node1306_r & ~pixel[520];
      node1311 = node1310_l;
      node1312 = node1310_r;
      node1313_r = node1297_r & pixel[440];
      node1313_l = node1297_r & ~pixel[440];
      node1314_r = node1313_l & pixel[387];
      node1314_l = node1313_l & ~pixel[387];
      node1315_r = node1314_l & pixel[543];
      node1315_l = node1314_l & ~pixel[543];
      node1316 = node1315_l;
      node1317 = node1315_r;
      node1318_r = node1314_r & pixel[546];
      node1318_l = node1314_r & ~pixel[546];
      node1319 = node1318_l;
      node1320 = node1318_r;
      node1321_r = node1313_r & pixel[610];
      node1321_l = node1313_r & ~pixel[610];
      node1322_r = node1321_l & pixel[525];
      node1322_l = node1321_l & ~pixel[525];
      node1323 = node1322_l;
      node1324 = node1322_r;
      node1325 = node1321_r;
      node1326_r = node1296_r & pixel[575];
      node1326_l = node1296_r & ~pixel[575];
      node1327_r = node1326_l & pixel[491];
      node1327_l = node1326_l & ~pixel[491];
      node1328_r = node1327_l & pixel[184];
      node1328_l = node1327_l & ~pixel[184];
      node1329_r = node1328_l & pixel[294];
      node1329_l = node1328_l & ~pixel[294];
      node1330 = node1329_l;
      node1331 = node1329_r;
      node1332_r = node1328_r & pixel[354];
      node1332_l = node1328_r & ~pixel[354];
      node1333 = node1332_l;
      node1334 = node1332_r;
      node1335_r = node1327_r & pixel[606];
      node1335_l = node1327_r & ~pixel[606];
      node1336_r = node1335_l & pixel[248];
      node1336_l = node1335_l & ~pixel[248];
      node1337 = node1336_l;
      node1338 = node1336_r;
      node1339_r = node1335_r & pixel[378];
      node1339_l = node1335_r & ~pixel[378];
      node1340 = node1339_l;
      node1341 = node1339_r;
      node1342_r = node1326_r & pixel[500];
      node1342_l = node1326_r & ~pixel[500];
      node1343_r = node1342_l & pixel[235];
      node1343_l = node1342_l & ~pixel[235];
      node1344_r = node1343_l & pixel[105];
      node1344_l = node1343_l & ~pixel[105];
      node1345 = node1344_l;
      node1346 = node1344_r;
      node1347_r = node1343_r & pixel[385];
      node1347_l = node1343_r & ~pixel[385];
      node1348 = node1347_l;
      node1349 = node1347_r;
      node1350_r = node1342_r & pixel[399];
      node1350_l = node1342_r & ~pixel[399];
      node1351_r = node1350_l & pixel[622];
      node1351_l = node1350_l & ~pixel[622];
      node1352 = node1351_l;
      node1353 = node1351_r;
      node1354_r = node1350_r & pixel[268];
      node1354_l = node1350_r & ~pixel[268];
      node1355 = node1354_l;
      node1356 = node1354_r;
      node1357_r = node1295_r & pixel[655];
      node1357_l = node1295_r & ~pixel[655];
      node1358_r = node1357_l & pixel[218];
      node1358_l = node1357_l & ~pixel[218];
      node1359_r = node1358_l & pixel[687];
      node1359_l = node1358_l & ~pixel[687];
      node1360_r = node1359_l & pixel[522];
      node1360_l = node1359_l & ~pixel[522];
      node1361_r = node1360_l & pixel[125];
      node1361_l = node1360_l & ~pixel[125];
      node1362 = node1361_l;
      node1363 = node1361_r;
      node1364_r = node1360_r & pixel[154];
      node1364_l = node1360_r & ~pixel[154];
      node1365 = node1364_l;
      node1366 = node1364_r;
      node1367 = node1359_r;
      node1368_r = node1358_r & pixel[269];
      node1368_l = node1358_r & ~pixel[269];
      node1369_r = node1368_l & pixel[401];
      node1369_l = node1368_l & ~pixel[401];
      node1370_r = node1369_l & pixel[262];
      node1370_l = node1369_l & ~pixel[262];
      node1371 = node1370_l;
      node1372 = node1370_r;
      node1373_r = node1369_r & pixel[567];
      node1373_l = node1369_r & ~pixel[567];
      node1374 = node1373_l;
      node1375 = node1373_r;
      node1376_r = node1368_r & pixel[159];
      node1376_l = node1368_r & ~pixel[159];
      node1377_r = node1376_l & pixel[381];
      node1377_l = node1376_l & ~pixel[381];
      node1378 = node1377_l;
      node1379 = node1377_r;
      node1380_r = node1376_r & pixel[405];
      node1380_l = node1376_r & ~pixel[405];
      node1381 = node1380_l;
      node1382 = node1380_r;
      node1383_r = node1357_r & pixel[456];
      node1383_l = node1357_r & ~pixel[456];
      node1384_r = node1383_l & pixel[551];
      node1384_l = node1383_l & ~pixel[551];
      node1385_r = node1384_l & pixel[682];
      node1385_l = node1384_l & ~pixel[682];
      node1386_r = node1385_l & pixel[514];
      node1386_l = node1385_l & ~pixel[514];
      node1387 = node1386_l;
      node1388 = node1386_r;
      node1389_r = node1385_r & pixel[454];
      node1389_l = node1385_r & ~pixel[454];
      node1390 = node1389_l;
      node1391 = node1389_r;
      node1392_r = node1384_r & pixel[515];
      node1392_l = node1384_r & ~pixel[515];
      node1393_r = node1392_l & pixel[352];
      node1393_l = node1392_l & ~pixel[352];
      node1394 = node1393_l;
      node1395 = node1393_r;
      node1396_r = node1392_r & pixel[377];
      node1396_l = node1392_r & ~pixel[377];
      node1397 = node1396_l;
      node1398 = node1396_r;
      node1399_r = node1383_r & pixel[354];
      node1399_l = node1383_r & ~pixel[354];
      node1400_r = node1399_l & pixel[435];
      node1400_l = node1399_l & ~pixel[435];
      node1401_r = node1400_l & pixel[157];
      node1401_l = node1400_l & ~pixel[157];
      node1402 = node1401_l;
      node1403 = node1401_r;
      node1404_r = node1400_r & pixel[510];
      node1404_l = node1400_r & ~pixel[510];
      node1405 = node1404_l;
      node1406 = node1404_r;
      node1407_r = node1399_r & pixel[468];
      node1407_l = node1399_r & ~pixel[468];
      node1408_r = node1407_l & pixel[485];
      node1408_l = node1407_l & ~pixel[485];
      node1409 = node1408_l;
      node1410 = node1408_r;
      node1411_r = node1407_r & pixel[207];
      node1411_l = node1407_r & ~pixel[207];
      node1412 = node1411_l;
      node1413 = node1411_r;
      node1414_r = node1174_r & pixel[292];
      node1414_l = node1174_r & ~pixel[292];
      node1415_r = node1414_l & pixel[468];
      node1415_l = node1414_l & ~pixel[468];
      node1416_r = node1415_l & pixel[618];
      node1416_l = node1415_l & ~pixel[618];
      node1417_r = node1416_l & pixel[101];
      node1417_l = node1416_l & ~pixel[101];
      node1418_r = node1417_l & pixel[267];
      node1418_l = node1417_l & ~pixel[267];
      node1419_r = node1418_l & pixel[436];
      node1419_l = node1418_l & ~pixel[436];
      node1420_r = node1419_l & pixel[543];
      node1420_l = node1419_l & ~pixel[543];
      node1421 = node1420_l;
      node1422 = node1420_r;
      node1423_r = node1419_r & pixel[184];
      node1423_l = node1419_r & ~pixel[184];
      node1424 = node1423_l;
      node1425 = node1423_r;
      node1426 = node1418_r;
      node1427_r = node1417_r & pixel[349];
      node1427_l = node1417_r & ~pixel[349];
      node1428_r = node1427_l & pixel[199];
      node1428_l = node1427_l & ~pixel[199];
      node1429_r = node1428_l & pixel[342];
      node1429_l = node1428_l & ~pixel[342];
      node1430 = node1429_l;
      node1431 = node1429_r;
      node1432 = node1428_r;
      node1433_r = node1427_r & pixel[552];
      node1433_l = node1427_r & ~pixel[552];
      node1434_r = node1433_l & pixel[581];
      node1434_l = node1433_l & ~pixel[581];
      node1435 = node1434_l;
      node1436 = node1434_r;
      node1437_r = node1433_r & pixel[297];
      node1437_l = node1433_r & ~pixel[297];
      node1438 = node1437_l;
      node1439 = node1437_r;
      node1440_r = node1416_r & pixel[550];
      node1440_l = node1416_r & ~pixel[550];
      node1441 = node1440_l;
      node1442 = node1440_r;
      node1443_r = node1415_r & pixel[262];
      node1443_l = node1415_r & ~pixel[262];
      node1444_r = node1443_l & pixel[100];
      node1444_l = node1443_l & ~pixel[100];
      node1445_r = node1444_l & pixel[183];
      node1445_l = node1444_l & ~pixel[183];
      node1446 = node1445_l;
      node1447 = node1445_r;
      node1448_r = node1444_r & pixel[259];
      node1448_l = node1444_r & ~pixel[259];
      node1449_r = node1448_l & pixel[432];
      node1449_l = node1448_l & ~pixel[432];
      node1450_r = node1449_l & pixel[490];
      node1450_l = node1449_l & ~pixel[490];
      node1451 = node1450_l;
      node1452 = node1450_r;
      node1453 = node1449_r;
      node1454_r = node1448_r & pixel[379];
      node1454_l = node1448_r & ~pixel[379];
      node1455 = node1454_l;
      node1456 = node1454_r;
      node1457_r = node1443_r & pixel[289];
      node1457_l = node1443_r & ~pixel[289];
      node1458_r = node1457_l & pixel[161];
      node1458_l = node1457_l & ~pixel[161];
      node1459_r = node1458_l & pixel[583];
      node1459_l = node1458_l & ~pixel[583];
      node1460 = node1459_l;
      node1461 = node1459_r;
      node1462 = node1458_r;
      node1463_r = node1457_r & pixel[508];
      node1463_l = node1457_r & ~pixel[508];
      node1464_r = node1463_l & pixel[511];
      node1464_l = node1463_l & ~pixel[511];
      node1465 = node1464_l;
      node1466 = node1464_r;
      node1467 = node1463_r;
      node1468_r = node1414_r & pixel[243];
      node1468_l = node1414_r & ~pixel[243];
      node1469_r = node1468_l & pixel[439];
      node1469_l = node1468_l & ~pixel[439];
      node1470_r = node1469_l & pixel[356];
      node1470_l = node1469_l & ~pixel[356];
      node1471_r = node1470_l & pixel[553];
      node1471_l = node1470_l & ~pixel[553];
      node1472_r = node1471_l & pixel[298];
      node1472_l = node1471_l & ~pixel[298];
      node1473_r = node1472_l & pixel[466];
      node1473_l = node1472_l & ~pixel[466];
      node1474 = node1473_l;
      node1475 = node1473_r;
      node1476_r = node1472_r & pixel[470];
      node1476_l = node1472_r & ~pixel[470];
      node1477 = node1476_l;
      node1478 = node1476_r;
      node1479_r = node1471_r & pixel[622];
      node1479_l = node1471_r & ~pixel[622];
      node1480_r = node1479_l & pixel[105];
      node1480_l = node1479_l & ~pixel[105];
      node1481 = node1480_l;
      node1482 = node1480_r;
      node1483 = node1479_r;
      node1484_r = node1470_r & pixel[535];
      node1484_l = node1470_r & ~pixel[535];
      node1485 = node1484_l;
      node1486 = node1484_r;
      node1487_r = node1469_r & pixel[402];
      node1487_l = node1469_r & ~pixel[402];
      node1488_r = node1487_l & pixel[151];
      node1488_l = node1487_l & ~pixel[151];
      node1489_r = node1488_l & pixel[468];
      node1489_l = node1488_l & ~pixel[468];
      node1490_r = node1489_l & pixel[456];
      node1490_l = node1489_l & ~pixel[456];
      node1491 = node1490_l;
      node1492 = node1490_r;
      node1493 = node1489_r;
      node1494_r = node1488_r & pixel[408];
      node1494_l = node1488_r & ~pixel[408];
      node1495 = node1494_l;
      node1496_r = node1494_r & pixel[260];
      node1496_l = node1494_r & ~pixel[260];
      node1497 = node1496_l;
      node1498 = node1496_r;
      node1499 = node1487_r;
      node1500_r = node1468_r & pixel[374];
      node1500_l = node1468_r & ~pixel[374];
      node1501_r = node1500_l & pixel[291];
      node1501_l = node1500_l & ~pixel[291];
      node1502_r = node1501_l & pixel[495];
      node1502_l = node1501_l & ~pixel[495];
      node1503 = node1502_l;
      node1504 = node1502_r;
      node1505_r = node1501_r & pixel[518];
      node1505_l = node1501_r & ~pixel[518];
      node1506 = node1505_l;
      node1507_r = node1505_r & pixel[408];
      node1507_l = node1505_r & ~pixel[408];
      node1508_r = node1507_l & pixel[153];
      node1508_l = node1507_l & ~pixel[153];
      node1509 = node1508_l;
      node1510 = node1508_r;
      node1511 = node1507_r;
      node1512_r = node1500_r & pixel[299];
      node1512_l = node1500_r & ~pixel[299];
      node1513_r = node1512_l & pixel[325];
      node1513_l = node1512_l & ~pixel[325];
      node1514 = node1513_l;
      node1515 = node1513_r;
      node1516_r = node1512_r & pixel[514];
      node1516_l = node1512_r & ~pixel[514];
      node1517 = node1516_l;
      node1518_r = node1516_r & pixel[525];
      node1518_l = node1516_r & ~pixel[525];
      node1519_r = node1518_l & pixel[320];
      node1519_l = node1518_l & ~pixel[320];
      node1520 = node1519_l;
      node1521 = node1519_r;
      node1522 = node1518_r;
      result0 = node32 | node35 | node47 | node49 | node62 | node66 | node73 | node85 | node99 | node102 | node103 | node136 | node140 | node151 | node159 | node188 | node218 | node264 | node299 | node301 | node311 | node318 | node866 | node873 | node874 | node883 | node902 | node903 | node906 | node915 | node936 | node945 | node959 | node968 | node976 | node978 | node979 | node982 | node987 | node999 | node1004 | node1011 | node1012 | node1014 | node1021 | node1027 | node1031 | node1043 | node1044 | node1046 | node1047 | node1053 | node1062 | node1065 | node1067 | node1083 | node1090 | node1098 | node1102 | node1112 | node1116 | node1118 | node1119 | node1126 | node1133 | node1134 | node1146 | node1149 | node1161 | node1173 | node1209 | node1231 | node1287 | node1403 | node1412;
      result1 = node91 | node370 | node399 | node403 | node557 | node572 | node579 | node582 | node587 | node618 | node619 | node666 | node686 | node690 | node719 | node794 | node1183 | node1309 | node1424;
      result2 = node11 | node25 | node48 | node95 | node109 | node190 | node199 | node210 | node211 | node217 | node229 | node242 | node247 | node265 | node268 | node271 | node278 | node281 | node337 | node404 | node417 | node419 | node434 | node448 | node452 | node460 | node465 | node473 | node479 | node509 | node524 | node528 | node558 | node564 | node580 | node583 | node604 | node614 | node625 | node629 | node700 | node707 | node708 | node731 | node776 | node792 | node799 | node851 | node857 | node884 | node887 | node890 | node958 | node1000 | node1003 | node1006 | node1007 | node1022 | node1028 | node1030 | node1036 | node1051 | node1056 | node1074 | node1087 | node1095 | node1131 | node1159 | node1165 | node1172 | node1185 | node1186 | node1189 | node1193 | node1197 | node1198 | node1200 | node1208 | node1212 | node1215 | node1223 | node1227 | node1230 | node1238 | node1240 | node1247 | node1252 | node1255 | node1259 | node1263 | node1279 | node1304 | node1317 | node1319 | node1333 | node1337 | node1341 | node1352 | node1353 | node1356 | node1363 | node1381 | node1397 | node1422 | node1425 | node1430 | node1436 | node1438 | node1439 | node1442 | node1447 | node1452 | node1453 | node1455 | node1461 | node1462 | node1481 | node1483 | node1486 | node1492 | node1503 | node1510 | node1511 | node1520 | node1522;
      result3 = node18 | node46 | node84 | node100 | node118 | node121 | node149 | node163 | node164 | node167 | node171 | node173 | node183 | node194 | node196 | node198 | node226 | node230 | node243 | node246 | node307 | node319 | node322 | node328 | node335 | node336 | node339 | node353 | node358 | node391 | node497 | node515 | node516 | node590 | node597 | node607 | node635 | node636 | node639 | node646 | node651 | node704 | node712 | node716 | node736 | node744 | node751 | node760 | node761 | node763 | node767 | node770 | node782 | node785 | node806 | node807 | node809 | node828 | node845 | node859 | node860 | node871 | node880 | node912 | node918 | node919 | node921 | node922 | node933 | node948 | node953 | node954 | node1054 | node1073 | node1086 | node1094 | node1097 | node1103 | node1109 | node1141 | node1144 | node1158 | node1162 | node1170 | node1171 | node1192 | node1221 | node1253 | node1284 | node1286 | node1325 | node1395 | node1409 | node1432 | node1441 | node1456 | node1495 | node1504 | node1509 | node1517;
      result4 = node10 | node13 | node78 | node87 | node92 | node110 | node135 | node139 | node143 | node222 | node240 | node270 | node286 | node288 | node294 | node295 | node298 | node341 | node367 | node371 | node383 | node415 | node426 | node427 | node436 | node442 | node444 | node445 | node457 | node468 | node480 | node508 | node512 | node594 | node610 | node638 | node643 | node673 | node729 | node732 | node743 | node802 | node863 | node898 | node950 | node964 | node971 | node983 | node1019 | node1127 | node1166 | node1205 | node1206 | node1244 | node1248 | node1256 | node1260 | node1269 | node1271 | node1302 | node1330 | node1340 | node1348 | node1362 | node1367 | node1374 | node1421 | node1467 | node1478 | node1515;
      result5 = node34 | node65 | node70 | node106 | node117 | node132 | node152 | node155 | node158 | node174 | node181 | node184 | node197 | node223 | node232 | node248 | node256 | node321 | node325 | node347 | node348 | node368 | node374 | node382 | node386 | node389 | node433 | node441 | node461 | node464 | node467 | node491 | node493 | node494 | node505 | node506 | node553 | node562 | node621 | node735 | node771 | node827 | node831 | node834 | node835 | node837 | node842 | node849 | node856 | node872 | node881 | node895 | node905 | node911 | node914 | node926 | node927 | node929 | node947 | node952 | node997 | node1061 | node1071 | node1082 | node1108 | node1153 | node1154 | node1220 | node1237 | node1268 | node1283 | node1290 | node1294 | node1301 | node1308 | node1312 | node1338 | node1371 | node1378 | node1382 | node1387 | node1391 | node1394 | node1402 | node1405 | node1474;
      result6 = node14 | node23 | node26 | node74 | node79 | node88 | node94 | node124 | node133 | node180 | node187 | node191 | node289 | node302 | node352 | node377 | node385 | node396 | node397 | node400 | node407 | node420 | node449 | node451 | node472 | node482 | node521 | node522 | node554 | node555 | node561 | node563 | node595 | node611 | node650 | node653 | node661 | node676 | node680 | node687 | node698 | node701 | node747 | node750 | node753 | node830 | node838 | node843 | node846 | node850 | node867 | node888 | node891 | node896 | node899 | node944 | node961 | node969 | node970 | node986 | node988 | node996 | node1018 | node1037 | node1081 | node1089 | node1111 | node1115 | node1123 | node1124 | node1130 | node1155 | node1213 | node1228 | node1245 | node1278 | node1320 | node1323 | node1324 | node1331 | node1345 | node1346 | node1349 | node1355 | node1365 | node1366 | node1426 | node1431 | node1446 | node1451 | node1460 | node1466 | node1475 | node1477 | node1482 | node1485 | node1491 | node1493 | node1498 | node1499 | node1514 | node1521;
      result7 = node17 | node20 | node21 | node31 | node38 | node41 | node55 | node59 | node63 | node156 | node207 | node208 | node215 | node225 | node239 | node254 | node255 | node258 | node263 | node279 | node282 | node306 | node310 | node313 | node314 | node326 | node346 | node355 | node406 | node437 | node531 | node537 | node546 | node575 | node603 | node606 | node674 | node723 | node739 | node791 | node801 | node813 | node1034 | node1048;
      result8 = node128 | node142 | node166 | node340 | node350 | node357 | node378 | node411 | node412 | node414 | node429 | node430 | node475 | node476 | node483 | node525 | node529 | node536 | node539 | node540 | node543 | node544 | node547 | node573 | node588 | node591 | node598 | node622 | node628 | node642 | node654 | node657 | node658 | node660 | node667 | node670 | node682 | node683 | node689 | node705 | node713 | node715 | node722 | node754 | node764 | node775 | node778 | node779 | node783 | node786 | node795 | node798 | node810 | node814 | node816 | node817 | node864 | node930 | node934 | node937 | node984 | node1066 | node1069 | node1101 | node1140 | node1143 | node1148 | node1182 | node1190 | node1241 | node1262 | node1275 | node1291 | node1293 | node1305 | node1311 | node1316 | node1334 | node1372 | node1375 | node1379 | node1388 | node1390 | node1398 | node1406 | node1410 | node1413 | node1435 | node1465 | node1497 | node1506;
      result9 = node39 | node42 | node56 | node58 | node71 | node77 | node107 | node120 | node125 | node127 | node148 | node170 | node214 | node233 | node237 | node259 | node266 | node285 | node293 | node329 | node375 | node390 | node458 | node490 | node498 | node500 | node501 | node513 | node532 | node576 | node613 | node626 | node645 | node669 | node677 | node697 | node720 | node728 | node738 | node746 | node768 | node963 | node1015 | node1035 | node1057 | node1199 | node1216 | node1224 | node1272 | node1276;

      tree_4 = {result9, result8, result7, result6, result5, result4, result3, result2, result1, result0};
    end
  endfunction

  function [9:0] tree_5;
    input [783:0] pixel;

    reg node0_r;
    reg node0_l;
    reg node1_r;
    reg node1_l;
    reg node2_r;
    reg node2_l;
    reg node3_r;
    reg node3_l;
    reg node4_r;
    reg node4_l;
    reg node5_r;
    reg node5_l;
    reg node6_r;
    reg node6_l;
    reg node7_r;
    reg node7_l;
    reg node8_r;
    reg node8_l;
    reg node9_r;
    reg node9_l;
    reg node10;
    reg node11;
    reg node12_r;
    reg node12_l;
    reg node13;
    reg node14;
    reg node15_r;
    reg node15_l;
    reg node16_r;
    reg node16_l;
    reg node17;
    reg node18;
    reg node19_r;
    reg node19_l;
    reg node20;
    reg node21;
    reg node22_r;
    reg node22_l;
    reg node23_r;
    reg node23_l;
    reg node24_r;
    reg node24_l;
    reg node25;
    reg node26;
    reg node27_r;
    reg node27_l;
    reg node28;
    reg node29;
    reg node30_r;
    reg node30_l;
    reg node31_r;
    reg node31_l;
    reg node32;
    reg node33;
    reg node34_r;
    reg node34_l;
    reg node35;
    reg node36;
    reg node37_r;
    reg node37_l;
    reg node38_r;
    reg node38_l;
    reg node39_r;
    reg node39_l;
    reg node40_r;
    reg node40_l;
    reg node41;
    reg node42;
    reg node43_r;
    reg node43_l;
    reg node44;
    reg node45;
    reg node46_r;
    reg node46_l;
    reg node47_r;
    reg node47_l;
    reg node48;
    reg node49;
    reg node50_r;
    reg node50_l;
    reg node51;
    reg node52;
    reg node53_r;
    reg node53_l;
    reg node54_r;
    reg node54_l;
    reg node55_r;
    reg node55_l;
    reg node56;
    reg node57;
    reg node58;
    reg node59_r;
    reg node59_l;
    reg node60;
    reg node61_r;
    reg node61_l;
    reg node62;
    reg node63;
    reg node64_r;
    reg node64_l;
    reg node65_r;
    reg node65_l;
    reg node66_r;
    reg node66_l;
    reg node67_r;
    reg node67_l;
    reg node68_r;
    reg node68_l;
    reg node69;
    reg node70;
    reg node71;
    reg node72_r;
    reg node72_l;
    reg node73_r;
    reg node73_l;
    reg node74;
    reg node75;
    reg node76_r;
    reg node76_l;
    reg node77;
    reg node78;
    reg node79_r;
    reg node79_l;
    reg node80_r;
    reg node80_l;
    reg node81_r;
    reg node81_l;
    reg node82;
    reg node83;
    reg node84_r;
    reg node84_l;
    reg node85;
    reg node86;
    reg node87_r;
    reg node87_l;
    reg node88_r;
    reg node88_l;
    reg node89;
    reg node90;
    reg node91;
    reg node92_r;
    reg node92_l;
    reg node93_r;
    reg node93_l;
    reg node94_r;
    reg node94_l;
    reg node95_r;
    reg node95_l;
    reg node96;
    reg node97;
    reg node98;
    reg node99_r;
    reg node99_l;
    reg node100_r;
    reg node100_l;
    reg node101;
    reg node102;
    reg node103_r;
    reg node103_l;
    reg node104;
    reg node105;
    reg node106_r;
    reg node106_l;
    reg node107_r;
    reg node107_l;
    reg node108_r;
    reg node108_l;
    reg node109;
    reg node110;
    reg node111_r;
    reg node111_l;
    reg node112;
    reg node113;
    reg node114_r;
    reg node114_l;
    reg node115_r;
    reg node115_l;
    reg node116;
    reg node117;
    reg node118;
    reg node119_r;
    reg node119_l;
    reg node120_r;
    reg node120_l;
    reg node121_r;
    reg node121_l;
    reg node122_r;
    reg node122_l;
    reg node123_r;
    reg node123_l;
    reg node124_r;
    reg node124_l;
    reg node125;
    reg node126;
    reg node127;
    reg node128_r;
    reg node128_l;
    reg node129;
    reg node130_r;
    reg node130_l;
    reg node131;
    reg node132;
    reg node133_r;
    reg node133_l;
    reg node134_r;
    reg node134_l;
    reg node135_r;
    reg node135_l;
    reg node136;
    reg node137;
    reg node138_r;
    reg node138_l;
    reg node139;
    reg node140;
    reg node141_r;
    reg node141_l;
    reg node142_r;
    reg node142_l;
    reg node143;
    reg node144;
    reg node145_r;
    reg node145_l;
    reg node146;
    reg node147;
    reg node148_r;
    reg node148_l;
    reg node149_r;
    reg node149_l;
    reg node150_r;
    reg node150_l;
    reg node151_r;
    reg node151_l;
    reg node152;
    reg node153;
    reg node154;
    reg node155_r;
    reg node155_l;
    reg node156_r;
    reg node156_l;
    reg node157;
    reg node158;
    reg node159_r;
    reg node159_l;
    reg node160;
    reg node161;
    reg node162_r;
    reg node162_l;
    reg node163_r;
    reg node163_l;
    reg node164;
    reg node165_r;
    reg node165_l;
    reg node166;
    reg node167;
    reg node168;
    reg node169_r;
    reg node169_l;
    reg node170_r;
    reg node170_l;
    reg node171_r;
    reg node171_l;
    reg node172_r;
    reg node172_l;
    reg node173_r;
    reg node173_l;
    reg node174;
    reg node175;
    reg node176_r;
    reg node176_l;
    reg node177;
    reg node178;
    reg node179_r;
    reg node179_l;
    reg node180_r;
    reg node180_l;
    reg node181;
    reg node182;
    reg node183_r;
    reg node183_l;
    reg node184;
    reg node185;
    reg node186_r;
    reg node186_l;
    reg node187_r;
    reg node187_l;
    reg node188_r;
    reg node188_l;
    reg node189;
    reg node190;
    reg node191;
    reg node192;
    reg node193_r;
    reg node193_l;
    reg node194_r;
    reg node194_l;
    reg node195_r;
    reg node195_l;
    reg node196_r;
    reg node196_l;
    reg node197;
    reg node198;
    reg node199_r;
    reg node199_l;
    reg node200;
    reg node201;
    reg node202_r;
    reg node202_l;
    reg node203;
    reg node204_r;
    reg node204_l;
    reg node205;
    reg node206;
    reg node207_r;
    reg node207_l;
    reg node208_r;
    reg node208_l;
    reg node209_r;
    reg node209_l;
    reg node210;
    reg node211;
    reg node212_r;
    reg node212_l;
    reg node213;
    reg node214;
    reg node215_r;
    reg node215_l;
    reg node216;
    reg node217;
    reg node218_r;
    reg node218_l;
    reg node219_r;
    reg node219_l;
    reg node220_r;
    reg node220_l;
    reg node221_r;
    reg node221_l;
    reg node222_r;
    reg node222_l;
    reg node223_r;
    reg node223_l;
    reg node224_r;
    reg node224_l;
    reg node225;
    reg node226;
    reg node227_r;
    reg node227_l;
    reg node228;
    reg node229;
    reg node230_r;
    reg node230_l;
    reg node231_r;
    reg node231_l;
    reg node232;
    reg node233;
    reg node234_r;
    reg node234_l;
    reg node235;
    reg node236;
    reg node237_r;
    reg node237_l;
    reg node238_r;
    reg node238_l;
    reg node239_r;
    reg node239_l;
    reg node240;
    reg node241;
    reg node242_r;
    reg node242_l;
    reg node243;
    reg node244;
    reg node245_r;
    reg node245_l;
    reg node246_r;
    reg node246_l;
    reg node247;
    reg node248;
    reg node249;
    reg node250_r;
    reg node250_l;
    reg node251_r;
    reg node251_l;
    reg node252_r;
    reg node252_l;
    reg node253_r;
    reg node253_l;
    reg node254;
    reg node255;
    reg node256_r;
    reg node256_l;
    reg node257;
    reg node258;
    reg node259_r;
    reg node259_l;
    reg node260_r;
    reg node260_l;
    reg node261;
    reg node262;
    reg node263_r;
    reg node263_l;
    reg node264;
    reg node265;
    reg node266_r;
    reg node266_l;
    reg node267_r;
    reg node267_l;
    reg node268_r;
    reg node268_l;
    reg node269;
    reg node270;
    reg node271_r;
    reg node271_l;
    reg node272;
    reg node273;
    reg node274_r;
    reg node274_l;
    reg node275_r;
    reg node275_l;
    reg node276;
    reg node277;
    reg node278;
    reg node279_r;
    reg node279_l;
    reg node280_r;
    reg node280_l;
    reg node281_r;
    reg node281_l;
    reg node282_r;
    reg node282_l;
    reg node283_r;
    reg node283_l;
    reg node284;
    reg node285;
    reg node286_r;
    reg node286_l;
    reg node287;
    reg node288;
    reg node289_r;
    reg node289_l;
    reg node290_r;
    reg node290_l;
    reg node291;
    reg node292;
    reg node293_r;
    reg node293_l;
    reg node294;
    reg node295;
    reg node296_r;
    reg node296_l;
    reg node297_r;
    reg node297_l;
    reg node298_r;
    reg node298_l;
    reg node299;
    reg node300;
    reg node301_r;
    reg node301_l;
    reg node302;
    reg node303;
    reg node304_r;
    reg node304_l;
    reg node305;
    reg node306_r;
    reg node306_l;
    reg node307;
    reg node308;
    reg node309_r;
    reg node309_l;
    reg node310_r;
    reg node310_l;
    reg node311_r;
    reg node311_l;
    reg node312_r;
    reg node312_l;
    reg node313;
    reg node314;
    reg node315_r;
    reg node315_l;
    reg node316;
    reg node317;
    reg node318_r;
    reg node318_l;
    reg node319_r;
    reg node319_l;
    reg node320;
    reg node321;
    reg node322_r;
    reg node322_l;
    reg node323;
    reg node324;
    reg node325_r;
    reg node325_l;
    reg node326_r;
    reg node326_l;
    reg node327_r;
    reg node327_l;
    reg node328;
    reg node329;
    reg node330_r;
    reg node330_l;
    reg node331;
    reg node332;
    reg node333_r;
    reg node333_l;
    reg node334_r;
    reg node334_l;
    reg node335;
    reg node336;
    reg node337_r;
    reg node337_l;
    reg node338;
    reg node339;
    reg node340_r;
    reg node340_l;
    reg node341_r;
    reg node341_l;
    reg node342_r;
    reg node342_l;
    reg node343_r;
    reg node343_l;
    reg node344_r;
    reg node344_l;
    reg node345_r;
    reg node345_l;
    reg node346;
    reg node347;
    reg node348_r;
    reg node348_l;
    reg node349;
    reg node350;
    reg node351_r;
    reg node351_l;
    reg node352_r;
    reg node352_l;
    reg node353;
    reg node354;
    reg node355_r;
    reg node355_l;
    reg node356;
    reg node357;
    reg node358_r;
    reg node358_l;
    reg node359_r;
    reg node359_l;
    reg node360_r;
    reg node360_l;
    reg node361;
    reg node362;
    reg node363_r;
    reg node363_l;
    reg node364;
    reg node365;
    reg node366_r;
    reg node366_l;
    reg node367_r;
    reg node367_l;
    reg node368;
    reg node369;
    reg node370_r;
    reg node370_l;
    reg node371;
    reg node372;
    reg node373_r;
    reg node373_l;
    reg node374_r;
    reg node374_l;
    reg node375_r;
    reg node375_l;
    reg node376_r;
    reg node376_l;
    reg node377;
    reg node378;
    reg node379_r;
    reg node379_l;
    reg node380;
    reg node381;
    reg node382_r;
    reg node382_l;
    reg node383_r;
    reg node383_l;
    reg node384;
    reg node385;
    reg node386_r;
    reg node386_l;
    reg node387;
    reg node388;
    reg node389_r;
    reg node389_l;
    reg node390_r;
    reg node390_l;
    reg node391_r;
    reg node391_l;
    reg node392;
    reg node393;
    reg node394_r;
    reg node394_l;
    reg node395;
    reg node396;
    reg node397;
    reg node398_r;
    reg node398_l;
    reg node399_r;
    reg node399_l;
    reg node400_r;
    reg node400_l;
    reg node401_r;
    reg node401_l;
    reg node402_r;
    reg node402_l;
    reg node403;
    reg node404;
    reg node405_r;
    reg node405_l;
    reg node406;
    reg node407;
    reg node408_r;
    reg node408_l;
    reg node409;
    reg node410;
    reg node411_r;
    reg node411_l;
    reg node412_r;
    reg node412_l;
    reg node413_r;
    reg node413_l;
    reg node414;
    reg node415;
    reg node416_r;
    reg node416_l;
    reg node417;
    reg node418;
    reg node419;
    reg node420_r;
    reg node420_l;
    reg node421_r;
    reg node421_l;
    reg node422_r;
    reg node422_l;
    reg node423_r;
    reg node423_l;
    reg node424;
    reg node425;
    reg node426;
    reg node427_r;
    reg node427_l;
    reg node428_r;
    reg node428_l;
    reg node429;
    reg node430;
    reg node431_r;
    reg node431_l;
    reg node432;
    reg node433;
    reg node434_r;
    reg node434_l;
    reg node435_r;
    reg node435_l;
    reg node436_r;
    reg node436_l;
    reg node437;
    reg node438;
    reg node439;
    reg node440_r;
    reg node440_l;
    reg node441_r;
    reg node441_l;
    reg node442;
    reg node443;
    reg node444_r;
    reg node444_l;
    reg node445;
    reg node446;
    reg node447_r;
    reg node447_l;
    reg node448_r;
    reg node448_l;
    reg node449_r;
    reg node449_l;
    reg node450_r;
    reg node450_l;
    reg node451_r;
    reg node451_l;
    reg node452_r;
    reg node452_l;
    reg node453_r;
    reg node453_l;
    reg node454_r;
    reg node454_l;
    reg node455;
    reg node456;
    reg node457_r;
    reg node457_l;
    reg node458;
    reg node459;
    reg node460_r;
    reg node460_l;
    reg node461_r;
    reg node461_l;
    reg node462;
    reg node463;
    reg node464_r;
    reg node464_l;
    reg node465;
    reg node466;
    reg node467_r;
    reg node467_l;
    reg node468_r;
    reg node468_l;
    reg node469_r;
    reg node469_l;
    reg node470;
    reg node471;
    reg node472_r;
    reg node472_l;
    reg node473;
    reg node474;
    reg node475_r;
    reg node475_l;
    reg node476_r;
    reg node476_l;
    reg node477;
    reg node478;
    reg node479_r;
    reg node479_l;
    reg node480;
    reg node481;
    reg node482_r;
    reg node482_l;
    reg node483_r;
    reg node483_l;
    reg node484_r;
    reg node484_l;
    reg node485_r;
    reg node485_l;
    reg node486;
    reg node487;
    reg node488_r;
    reg node488_l;
    reg node489;
    reg node490;
    reg node491_r;
    reg node491_l;
    reg node492_r;
    reg node492_l;
    reg node493;
    reg node494;
    reg node495_r;
    reg node495_l;
    reg node496;
    reg node497;
    reg node498_r;
    reg node498_l;
    reg node499_r;
    reg node499_l;
    reg node500_r;
    reg node500_l;
    reg node501;
    reg node502;
    reg node503_r;
    reg node503_l;
    reg node504;
    reg node505;
    reg node506_r;
    reg node506_l;
    reg node507_r;
    reg node507_l;
    reg node508;
    reg node509;
    reg node510;
    reg node511_r;
    reg node511_l;
    reg node512_r;
    reg node512_l;
    reg node513_r;
    reg node513_l;
    reg node514_r;
    reg node514_l;
    reg node515;
    reg node516_r;
    reg node516_l;
    reg node517;
    reg node518;
    reg node519_r;
    reg node519_l;
    reg node520_r;
    reg node520_l;
    reg node521;
    reg node522;
    reg node523;
    reg node524_r;
    reg node524_l;
    reg node525_r;
    reg node525_l;
    reg node526_r;
    reg node526_l;
    reg node527;
    reg node528;
    reg node529_r;
    reg node529_l;
    reg node530;
    reg node531;
    reg node532;
    reg node533_r;
    reg node533_l;
    reg node534_r;
    reg node534_l;
    reg node535_r;
    reg node535_l;
    reg node536_r;
    reg node536_l;
    reg node537;
    reg node538;
    reg node539;
    reg node540_r;
    reg node540_l;
    reg node541_r;
    reg node541_l;
    reg node542;
    reg node543;
    reg node544;
    reg node545_r;
    reg node545_l;
    reg node546_r;
    reg node546_l;
    reg node547_r;
    reg node547_l;
    reg node548;
    reg node549;
    reg node550_r;
    reg node550_l;
    reg node551;
    reg node552;
    reg node553_r;
    reg node553_l;
    reg node554_r;
    reg node554_l;
    reg node555;
    reg node556;
    reg node557_r;
    reg node557_l;
    reg node558;
    reg node559;
    reg node560_r;
    reg node560_l;
    reg node561_r;
    reg node561_l;
    reg node562_r;
    reg node562_l;
    reg node563_r;
    reg node563_l;
    reg node564_r;
    reg node564_l;
    reg node565_r;
    reg node565_l;
    reg node566;
    reg node567;
    reg node568_r;
    reg node568_l;
    reg node569;
    reg node570;
    reg node571_r;
    reg node571_l;
    reg node572_r;
    reg node572_l;
    reg node573;
    reg node574;
    reg node575_r;
    reg node575_l;
    reg node576;
    reg node577;
    reg node578_r;
    reg node578_l;
    reg node579_r;
    reg node579_l;
    reg node580_r;
    reg node580_l;
    reg node581;
    reg node582;
    reg node583_r;
    reg node583_l;
    reg node584;
    reg node585;
    reg node586_r;
    reg node586_l;
    reg node587_r;
    reg node587_l;
    reg node588;
    reg node589;
    reg node590_r;
    reg node590_l;
    reg node591;
    reg node592;
    reg node593_r;
    reg node593_l;
    reg node594_r;
    reg node594_l;
    reg node595_r;
    reg node595_l;
    reg node596_r;
    reg node596_l;
    reg node597;
    reg node598;
    reg node599_r;
    reg node599_l;
    reg node600;
    reg node601;
    reg node602_r;
    reg node602_l;
    reg node603_r;
    reg node603_l;
    reg node604;
    reg node605;
    reg node606_r;
    reg node606_l;
    reg node607;
    reg node608;
    reg node609_r;
    reg node609_l;
    reg node610_r;
    reg node610_l;
    reg node611_r;
    reg node611_l;
    reg node612;
    reg node613;
    reg node614_r;
    reg node614_l;
    reg node615;
    reg node616;
    reg node617_r;
    reg node617_l;
    reg node618_r;
    reg node618_l;
    reg node619;
    reg node620;
    reg node621_r;
    reg node621_l;
    reg node622;
    reg node623;
    reg node624_r;
    reg node624_l;
    reg node625_r;
    reg node625_l;
    reg node626_r;
    reg node626_l;
    reg node627_r;
    reg node627_l;
    reg node628_r;
    reg node628_l;
    reg node629;
    reg node630;
    reg node631_r;
    reg node631_l;
    reg node632;
    reg node633;
    reg node634_r;
    reg node634_l;
    reg node635_r;
    reg node635_l;
    reg node636;
    reg node637;
    reg node638_r;
    reg node638_l;
    reg node639;
    reg node640;
    reg node641_r;
    reg node641_l;
    reg node642_r;
    reg node642_l;
    reg node643_r;
    reg node643_l;
    reg node644;
    reg node645;
    reg node646_r;
    reg node646_l;
    reg node647;
    reg node648;
    reg node649_r;
    reg node649_l;
    reg node650_r;
    reg node650_l;
    reg node651;
    reg node652;
    reg node653_r;
    reg node653_l;
    reg node654;
    reg node655;
    reg node656_r;
    reg node656_l;
    reg node657_r;
    reg node657_l;
    reg node658_r;
    reg node658_l;
    reg node659_r;
    reg node659_l;
    reg node660;
    reg node661;
    reg node662;
    reg node663_r;
    reg node663_l;
    reg node664_r;
    reg node664_l;
    reg node665;
    reg node666;
    reg node667_r;
    reg node667_l;
    reg node668;
    reg node669;
    reg node670_r;
    reg node670_l;
    reg node671_r;
    reg node671_l;
    reg node672_r;
    reg node672_l;
    reg node673;
    reg node674;
    reg node675_r;
    reg node675_l;
    reg node676;
    reg node677;
    reg node678_r;
    reg node678_l;
    reg node679_r;
    reg node679_l;
    reg node680;
    reg node681;
    reg node682_r;
    reg node682_l;
    reg node683;
    reg node684;
    reg node685_r;
    reg node685_l;
    reg node686_r;
    reg node686_l;
    reg node687_r;
    reg node687_l;
    reg node688_r;
    reg node688_l;
    reg node689_r;
    reg node689_l;
    reg node690_r;
    reg node690_l;
    reg node691_r;
    reg node691_l;
    reg node692;
    reg node693;
    reg node694_r;
    reg node694_l;
    reg node695;
    reg node696;
    reg node697_r;
    reg node697_l;
    reg node698_r;
    reg node698_l;
    reg node699;
    reg node700;
    reg node701_r;
    reg node701_l;
    reg node702;
    reg node703;
    reg node704_r;
    reg node704_l;
    reg node705_r;
    reg node705_l;
    reg node706_r;
    reg node706_l;
    reg node707;
    reg node708;
    reg node709_r;
    reg node709_l;
    reg node710;
    reg node711;
    reg node712_r;
    reg node712_l;
    reg node713_r;
    reg node713_l;
    reg node714;
    reg node715;
    reg node716_r;
    reg node716_l;
    reg node717;
    reg node718;
    reg node719_r;
    reg node719_l;
    reg node720_r;
    reg node720_l;
    reg node721_r;
    reg node721_l;
    reg node722_r;
    reg node722_l;
    reg node723;
    reg node724;
    reg node725_r;
    reg node725_l;
    reg node726;
    reg node727;
    reg node728_r;
    reg node728_l;
    reg node729_r;
    reg node729_l;
    reg node730;
    reg node731;
    reg node732_r;
    reg node732_l;
    reg node733;
    reg node734;
    reg node735_r;
    reg node735_l;
    reg node736_r;
    reg node736_l;
    reg node737;
    reg node738;
    reg node739_r;
    reg node739_l;
    reg node740_r;
    reg node740_l;
    reg node741;
    reg node742;
    reg node743_r;
    reg node743_l;
    reg node744;
    reg node745;
    reg node746_r;
    reg node746_l;
    reg node747_r;
    reg node747_l;
    reg node748_r;
    reg node748_l;
    reg node749_r;
    reg node749_l;
    reg node750_r;
    reg node750_l;
    reg node751;
    reg node752;
    reg node753_r;
    reg node753_l;
    reg node754;
    reg node755;
    reg node756_r;
    reg node756_l;
    reg node757_r;
    reg node757_l;
    reg node758;
    reg node759;
    reg node760_r;
    reg node760_l;
    reg node761;
    reg node762;
    reg node763_r;
    reg node763_l;
    reg node764_r;
    reg node764_l;
    reg node765_r;
    reg node765_l;
    reg node766;
    reg node767;
    reg node768;
    reg node769_r;
    reg node769_l;
    reg node770_r;
    reg node770_l;
    reg node771;
    reg node772;
    reg node773_r;
    reg node773_l;
    reg node774;
    reg node775;
    reg node776_r;
    reg node776_l;
    reg node777_r;
    reg node777_l;
    reg node778_r;
    reg node778_l;
    reg node779_r;
    reg node779_l;
    reg node780;
    reg node781;
    reg node782_r;
    reg node782_l;
    reg node783;
    reg node784;
    reg node785_r;
    reg node785_l;
    reg node786_r;
    reg node786_l;
    reg node787;
    reg node788;
    reg node789_r;
    reg node789_l;
    reg node790;
    reg node791;
    reg node792_r;
    reg node792_l;
    reg node793_r;
    reg node793_l;
    reg node794_r;
    reg node794_l;
    reg node795;
    reg node796;
    reg node797_r;
    reg node797_l;
    reg node798;
    reg node799;
    reg node800_r;
    reg node800_l;
    reg node801_r;
    reg node801_l;
    reg node802;
    reg node803;
    reg node804_r;
    reg node804_l;
    reg node805;
    reg node806;
    reg node807_r;
    reg node807_l;
    reg node808_r;
    reg node808_l;
    reg node809_r;
    reg node809_l;
    reg node810_r;
    reg node810_l;
    reg node811_r;
    reg node811_l;
    reg node812_r;
    reg node812_l;
    reg node813;
    reg node814;
    reg node815_r;
    reg node815_l;
    reg node816;
    reg node817;
    reg node818_r;
    reg node818_l;
    reg node819_r;
    reg node819_l;
    reg node820;
    reg node821;
    reg node822_r;
    reg node822_l;
    reg node823;
    reg node824;
    reg node825_r;
    reg node825_l;
    reg node826_r;
    reg node826_l;
    reg node827_r;
    reg node827_l;
    reg node828;
    reg node829;
    reg node830_r;
    reg node830_l;
    reg node831;
    reg node832;
    reg node833;
    reg node834_r;
    reg node834_l;
    reg node835_r;
    reg node835_l;
    reg node836;
    reg node837;
    reg node838_r;
    reg node838_l;
    reg node839_r;
    reg node839_l;
    reg node840;
    reg node841;
    reg node842_r;
    reg node842_l;
    reg node843;
    reg node844_r;
    reg node844_l;
    reg node845;
    reg node846;
    reg node847_r;
    reg node847_l;
    reg node848_r;
    reg node848_l;
    reg node849_r;
    reg node849_l;
    reg node850_r;
    reg node850_l;
    reg node851_r;
    reg node851_l;
    reg node852;
    reg node853;
    reg node854_r;
    reg node854_l;
    reg node855;
    reg node856;
    reg node857_r;
    reg node857_l;
    reg node858_r;
    reg node858_l;
    reg node859;
    reg node860;
    reg node861_r;
    reg node861_l;
    reg node862;
    reg node863;
    reg node864_r;
    reg node864_l;
    reg node865_r;
    reg node865_l;
    reg node866_r;
    reg node866_l;
    reg node867;
    reg node868;
    reg node869_r;
    reg node869_l;
    reg node870;
    reg node871;
    reg node872_r;
    reg node872_l;
    reg node873_r;
    reg node873_l;
    reg node874;
    reg node875;
    reg node876_r;
    reg node876_l;
    reg node877;
    reg node878;
    reg node879_r;
    reg node879_l;
    reg node880_r;
    reg node880_l;
    reg node881_r;
    reg node881_l;
    reg node882_r;
    reg node882_l;
    reg node883;
    reg node884;
    reg node885_r;
    reg node885_l;
    reg node886;
    reg node887;
    reg node888_r;
    reg node888_l;
    reg node889_r;
    reg node889_l;
    reg node890;
    reg node891;
    reg node892_r;
    reg node892_l;
    reg node893;
    reg node894;
    reg node895_r;
    reg node895_l;
    reg node896_r;
    reg node896_l;
    reg node897_r;
    reg node897_l;
    reg node898;
    reg node899;
    reg node900_r;
    reg node900_l;
    reg node901;
    reg node902;
    reg node903_r;
    reg node903_l;
    reg node904_r;
    reg node904_l;
    reg node905;
    reg node906;
    reg node907_r;
    reg node907_l;
    reg node908;
    reg node909;
    reg node910_r;
    reg node910_l;
    reg node911_r;
    reg node911_l;
    reg node912_r;
    reg node912_l;
    reg node913_r;
    reg node913_l;
    reg node914_r;
    reg node914_l;
    reg node915_r;
    reg node915_l;
    reg node916_r;
    reg node916_l;
    reg node917_r;
    reg node917_l;
    reg node918_r;
    reg node918_l;
    reg node919;
    reg node920;
    reg node921_r;
    reg node921_l;
    reg node922;
    reg node923;
    reg node924_r;
    reg node924_l;
    reg node925_r;
    reg node925_l;
    reg node926;
    reg node927;
    reg node928_r;
    reg node928_l;
    reg node929;
    reg node930;
    reg node931_r;
    reg node931_l;
    reg node932_r;
    reg node932_l;
    reg node933_r;
    reg node933_l;
    reg node934;
    reg node935;
    reg node936_r;
    reg node936_l;
    reg node937;
    reg node938;
    reg node939_r;
    reg node939_l;
    reg node940_r;
    reg node940_l;
    reg node941;
    reg node942;
    reg node943;
    reg node944_r;
    reg node944_l;
    reg node945_r;
    reg node945_l;
    reg node946_r;
    reg node946_l;
    reg node947_r;
    reg node947_l;
    reg node948;
    reg node949;
    reg node950_r;
    reg node950_l;
    reg node951;
    reg node952;
    reg node953_r;
    reg node953_l;
    reg node954_r;
    reg node954_l;
    reg node955;
    reg node956;
    reg node957_r;
    reg node957_l;
    reg node958;
    reg node959;
    reg node960_r;
    reg node960_l;
    reg node961_r;
    reg node961_l;
    reg node962_r;
    reg node962_l;
    reg node963;
    reg node964;
    reg node965;
    reg node966_r;
    reg node966_l;
    reg node967_r;
    reg node967_l;
    reg node968;
    reg node969;
    reg node970;
    reg node971_r;
    reg node971_l;
    reg node972_r;
    reg node972_l;
    reg node973_r;
    reg node973_l;
    reg node974_r;
    reg node974_l;
    reg node975_r;
    reg node975_l;
    reg node976;
    reg node977;
    reg node978_r;
    reg node978_l;
    reg node979;
    reg node980;
    reg node981_r;
    reg node981_l;
    reg node982_r;
    reg node982_l;
    reg node983;
    reg node984;
    reg node985_r;
    reg node985_l;
    reg node986;
    reg node987;
    reg node988_r;
    reg node988_l;
    reg node989_r;
    reg node989_l;
    reg node990_r;
    reg node990_l;
    reg node991;
    reg node992;
    reg node993_r;
    reg node993_l;
    reg node994;
    reg node995;
    reg node996_r;
    reg node996_l;
    reg node997_r;
    reg node997_l;
    reg node998;
    reg node999;
    reg node1000_r;
    reg node1000_l;
    reg node1001;
    reg node1002;
    reg node1003_r;
    reg node1003_l;
    reg node1004_r;
    reg node1004_l;
    reg node1005_r;
    reg node1005_l;
    reg node1006_r;
    reg node1006_l;
    reg node1007;
    reg node1008;
    reg node1009_r;
    reg node1009_l;
    reg node1010;
    reg node1011;
    reg node1012_r;
    reg node1012_l;
    reg node1013_r;
    reg node1013_l;
    reg node1014;
    reg node1015;
    reg node1016_r;
    reg node1016_l;
    reg node1017;
    reg node1018;
    reg node1019_r;
    reg node1019_l;
    reg node1020_r;
    reg node1020_l;
    reg node1021_r;
    reg node1021_l;
    reg node1022;
    reg node1023;
    reg node1024_r;
    reg node1024_l;
    reg node1025;
    reg node1026;
    reg node1027;
    reg node1028_r;
    reg node1028_l;
    reg node1029_r;
    reg node1029_l;
    reg node1030_r;
    reg node1030_l;
    reg node1031_r;
    reg node1031_l;
    reg node1032_r;
    reg node1032_l;
    reg node1033_r;
    reg node1033_l;
    reg node1034;
    reg node1035;
    reg node1036_r;
    reg node1036_l;
    reg node1037;
    reg node1038;
    reg node1039_r;
    reg node1039_l;
    reg node1040;
    reg node1041;
    reg node1042_r;
    reg node1042_l;
    reg node1043_r;
    reg node1043_l;
    reg node1044_r;
    reg node1044_l;
    reg node1045;
    reg node1046;
    reg node1047_r;
    reg node1047_l;
    reg node1048;
    reg node1049;
    reg node1050_r;
    reg node1050_l;
    reg node1051_r;
    reg node1051_l;
    reg node1052;
    reg node1053;
    reg node1054_r;
    reg node1054_l;
    reg node1055;
    reg node1056;
    reg node1057_r;
    reg node1057_l;
    reg node1058_r;
    reg node1058_l;
    reg node1059_r;
    reg node1059_l;
    reg node1060_r;
    reg node1060_l;
    reg node1061;
    reg node1062;
    reg node1063_r;
    reg node1063_l;
    reg node1064;
    reg node1065;
    reg node1066_r;
    reg node1066_l;
    reg node1067_r;
    reg node1067_l;
    reg node1068;
    reg node1069;
    reg node1070_r;
    reg node1070_l;
    reg node1071;
    reg node1072;
    reg node1073_r;
    reg node1073_l;
    reg node1074_r;
    reg node1074_l;
    reg node1075_r;
    reg node1075_l;
    reg node1076;
    reg node1077;
    reg node1078_r;
    reg node1078_l;
    reg node1079;
    reg node1080;
    reg node1081_r;
    reg node1081_l;
    reg node1082_r;
    reg node1082_l;
    reg node1083;
    reg node1084;
    reg node1085_r;
    reg node1085_l;
    reg node1086;
    reg node1087;
    reg node1088_r;
    reg node1088_l;
    reg node1089_r;
    reg node1089_l;
    reg node1090_r;
    reg node1090_l;
    reg node1091_r;
    reg node1091_l;
    reg node1092_r;
    reg node1092_l;
    reg node1093;
    reg node1094;
    reg node1095_r;
    reg node1095_l;
    reg node1096;
    reg node1097;
    reg node1098_r;
    reg node1098_l;
    reg node1099_r;
    reg node1099_l;
    reg node1100;
    reg node1101;
    reg node1102_r;
    reg node1102_l;
    reg node1103;
    reg node1104;
    reg node1105_r;
    reg node1105_l;
    reg node1106_r;
    reg node1106_l;
    reg node1107_r;
    reg node1107_l;
    reg node1108;
    reg node1109;
    reg node1110_r;
    reg node1110_l;
    reg node1111;
    reg node1112;
    reg node1113_r;
    reg node1113_l;
    reg node1114_r;
    reg node1114_l;
    reg node1115;
    reg node1116;
    reg node1117_r;
    reg node1117_l;
    reg node1118;
    reg node1119;
    reg node1120_r;
    reg node1120_l;
    reg node1121_r;
    reg node1121_l;
    reg node1122_r;
    reg node1122_l;
    reg node1123_r;
    reg node1123_l;
    reg node1124;
    reg node1125;
    reg node1126_r;
    reg node1126_l;
    reg node1127;
    reg node1128;
    reg node1129_r;
    reg node1129_l;
    reg node1130_r;
    reg node1130_l;
    reg node1131;
    reg node1132;
    reg node1133_r;
    reg node1133_l;
    reg node1134;
    reg node1135;
    reg node1136_r;
    reg node1136_l;
    reg node1137_r;
    reg node1137_l;
    reg node1138_r;
    reg node1138_l;
    reg node1139;
    reg node1140;
    reg node1141_r;
    reg node1141_l;
    reg node1142;
    reg node1143;
    reg node1144_r;
    reg node1144_l;
    reg node1145_r;
    reg node1145_l;
    reg node1146;
    reg node1147;
    reg node1148_r;
    reg node1148_l;
    reg node1149;
    reg node1150;
    reg node1151_r;
    reg node1151_l;
    reg node1152_r;
    reg node1152_l;
    reg node1153_r;
    reg node1153_l;
    reg node1154_r;
    reg node1154_l;
    reg node1155_r;
    reg node1155_l;
    reg node1156_r;
    reg node1156_l;
    reg node1157_r;
    reg node1157_l;
    reg node1158;
    reg node1159;
    reg node1160_r;
    reg node1160_l;
    reg node1161;
    reg node1162;
    reg node1163_r;
    reg node1163_l;
    reg node1164_r;
    reg node1164_l;
    reg node1165;
    reg node1166;
    reg node1167_r;
    reg node1167_l;
    reg node1168;
    reg node1169;
    reg node1170_r;
    reg node1170_l;
    reg node1171_r;
    reg node1171_l;
    reg node1172_r;
    reg node1172_l;
    reg node1173;
    reg node1174;
    reg node1175_r;
    reg node1175_l;
    reg node1176;
    reg node1177;
    reg node1178_r;
    reg node1178_l;
    reg node1179_r;
    reg node1179_l;
    reg node1180;
    reg node1181;
    reg node1182_r;
    reg node1182_l;
    reg node1183;
    reg node1184;
    reg node1185_r;
    reg node1185_l;
    reg node1186_r;
    reg node1186_l;
    reg node1187_r;
    reg node1187_l;
    reg node1188_r;
    reg node1188_l;
    reg node1189;
    reg node1190;
    reg node1191;
    reg node1192_r;
    reg node1192_l;
    reg node1193_r;
    reg node1193_l;
    reg node1194;
    reg node1195;
    reg node1196;
    reg node1197_r;
    reg node1197_l;
    reg node1198;
    reg node1199_r;
    reg node1199_l;
    reg node1200;
    reg node1201;
    reg node1202_r;
    reg node1202_l;
    reg node1203_r;
    reg node1203_l;
    reg node1204_r;
    reg node1204_l;
    reg node1205_r;
    reg node1205_l;
    reg node1206_r;
    reg node1206_l;
    reg node1207;
    reg node1208;
    reg node1209_r;
    reg node1209_l;
    reg node1210;
    reg node1211;
    reg node1212_r;
    reg node1212_l;
    reg node1213_r;
    reg node1213_l;
    reg node1214;
    reg node1215;
    reg node1216_r;
    reg node1216_l;
    reg node1217;
    reg node1218;
    reg node1219_r;
    reg node1219_l;
    reg node1220_r;
    reg node1220_l;
    reg node1221;
    reg node1222;
    reg node1223_r;
    reg node1223_l;
    reg node1224_r;
    reg node1224_l;
    reg node1225;
    reg node1226;
    reg node1227_r;
    reg node1227_l;
    reg node1228;
    reg node1229;
    reg node1230_r;
    reg node1230_l;
    reg node1231_r;
    reg node1231_l;
    reg node1232_r;
    reg node1232_l;
    reg node1233_r;
    reg node1233_l;
    reg node1234;
    reg node1235;
    reg node1236;
    reg node1237_r;
    reg node1237_l;
    reg node1238;
    reg node1239_r;
    reg node1239_l;
    reg node1240;
    reg node1241;
    reg node1242_r;
    reg node1242_l;
    reg node1243_r;
    reg node1243_l;
    reg node1244_r;
    reg node1244_l;
    reg node1245;
    reg node1246;
    reg node1247_r;
    reg node1247_l;
    reg node1248;
    reg node1249;
    reg node1250_r;
    reg node1250_l;
    reg node1251_r;
    reg node1251_l;
    reg node1252;
    reg node1253;
    reg node1254_r;
    reg node1254_l;
    reg node1255;
    reg node1256;
    reg node1257_r;
    reg node1257_l;
    reg node1258_r;
    reg node1258_l;
    reg node1259_r;
    reg node1259_l;
    reg node1260_r;
    reg node1260_l;
    reg node1261_r;
    reg node1261_l;
    reg node1262_r;
    reg node1262_l;
    reg node1263;
    reg node1264;
    reg node1265;
    reg node1266_r;
    reg node1266_l;
    reg node1267_r;
    reg node1267_l;
    reg node1268;
    reg node1269;
    reg node1270_r;
    reg node1270_l;
    reg node1271;
    reg node1272;
    reg node1273_r;
    reg node1273_l;
    reg node1274_r;
    reg node1274_l;
    reg node1275;
    reg node1276_r;
    reg node1276_l;
    reg node1277;
    reg node1278;
    reg node1279_r;
    reg node1279_l;
    reg node1280_r;
    reg node1280_l;
    reg node1281;
    reg node1282;
    reg node1283_r;
    reg node1283_l;
    reg node1284;
    reg node1285;
    reg node1286_r;
    reg node1286_l;
    reg node1287_r;
    reg node1287_l;
    reg node1288_r;
    reg node1288_l;
    reg node1289_r;
    reg node1289_l;
    reg node1290;
    reg node1291;
    reg node1292_r;
    reg node1292_l;
    reg node1293;
    reg node1294;
    reg node1295_r;
    reg node1295_l;
    reg node1296_r;
    reg node1296_l;
    reg node1297;
    reg node1298;
    reg node1299_r;
    reg node1299_l;
    reg node1300;
    reg node1301;
    reg node1302_r;
    reg node1302_l;
    reg node1303_r;
    reg node1303_l;
    reg node1304_r;
    reg node1304_l;
    reg node1305;
    reg node1306;
    reg node1307_r;
    reg node1307_l;
    reg node1308;
    reg node1309;
    reg node1310_r;
    reg node1310_l;
    reg node1311_r;
    reg node1311_l;
    reg node1312;
    reg node1313;
    reg node1314_r;
    reg node1314_l;
    reg node1315;
    reg node1316;
    reg node1317_r;
    reg node1317_l;
    reg node1318_r;
    reg node1318_l;
    reg node1319_r;
    reg node1319_l;
    reg node1320_r;
    reg node1320_l;
    reg node1321;
    reg node1322_r;
    reg node1322_l;
    reg node1323;
    reg node1324;
    reg node1325_r;
    reg node1325_l;
    reg node1326_r;
    reg node1326_l;
    reg node1327;
    reg node1328;
    reg node1329_r;
    reg node1329_l;
    reg node1330;
    reg node1331;
    reg node1332_r;
    reg node1332_l;
    reg node1333_r;
    reg node1333_l;
    reg node1334_r;
    reg node1334_l;
    reg node1335;
    reg node1336;
    reg node1337;
    reg node1338_r;
    reg node1338_l;
    reg node1339;
    reg node1340_r;
    reg node1340_l;
    reg node1341;
    reg node1342;
    reg node1343_r;
    reg node1343_l;
    reg node1344_r;
    reg node1344_l;
    reg node1345_r;
    reg node1345_l;
    reg node1346_r;
    reg node1346_l;
    reg node1347;
    reg node1348;
    reg node1349_r;
    reg node1349_l;
    reg node1350;
    reg node1351;
    reg node1352_r;
    reg node1352_l;
    reg node1353_r;
    reg node1353_l;
    reg node1354;
    reg node1355;
    reg node1356_r;
    reg node1356_l;
    reg node1357;
    reg node1358;
    reg node1359_r;
    reg node1359_l;
    reg node1360_r;
    reg node1360_l;
    reg node1361_r;
    reg node1361_l;
    reg node1362;
    reg node1363;
    reg node1364_r;
    reg node1364_l;
    reg node1365;
    reg node1366;
    reg node1367_r;
    reg node1367_l;
    reg node1368_r;
    reg node1368_l;
    reg node1369;
    reg node1370;
    reg node1371_r;
    reg node1371_l;
    reg node1372;
    reg node1373;
    reg node1374_r;
    reg node1374_l;
    reg node1375_r;
    reg node1375_l;
    reg node1376_r;
    reg node1376_l;
    reg node1377_r;
    reg node1377_l;
    reg node1378_r;
    reg node1378_l;
    reg node1379_r;
    reg node1379_l;
    reg node1380_r;
    reg node1380_l;
    reg node1381_r;
    reg node1381_l;
    reg node1382;
    reg node1383;
    reg node1384_r;
    reg node1384_l;
    reg node1385;
    reg node1386;
    reg node1387_r;
    reg node1387_l;
    reg node1388_r;
    reg node1388_l;
    reg node1389;
    reg node1390;
    reg node1391_r;
    reg node1391_l;
    reg node1392;
    reg node1393;
    reg node1394_r;
    reg node1394_l;
    reg node1395_r;
    reg node1395_l;
    reg node1396_r;
    reg node1396_l;
    reg node1397;
    reg node1398;
    reg node1399_r;
    reg node1399_l;
    reg node1400;
    reg node1401;
    reg node1402_r;
    reg node1402_l;
    reg node1403_r;
    reg node1403_l;
    reg node1404;
    reg node1405;
    reg node1406_r;
    reg node1406_l;
    reg node1407;
    reg node1408;
    reg node1409_r;
    reg node1409_l;
    reg node1410_r;
    reg node1410_l;
    reg node1411_r;
    reg node1411_l;
    reg node1412_r;
    reg node1412_l;
    reg node1413;
    reg node1414;
    reg node1415_r;
    reg node1415_l;
    reg node1416;
    reg node1417;
    reg node1418_r;
    reg node1418_l;
    reg node1419_r;
    reg node1419_l;
    reg node1420;
    reg node1421;
    reg node1422_r;
    reg node1422_l;
    reg node1423;
    reg node1424;
    reg node1425_r;
    reg node1425_l;
    reg node1426_r;
    reg node1426_l;
    reg node1427_r;
    reg node1427_l;
    reg node1428;
    reg node1429;
    reg node1430_r;
    reg node1430_l;
    reg node1431;
    reg node1432;
    reg node1433_r;
    reg node1433_l;
    reg node1434_r;
    reg node1434_l;
    reg node1435;
    reg node1436;
    reg node1437_r;
    reg node1437_l;
    reg node1438;
    reg node1439;
    reg node1440_r;
    reg node1440_l;
    reg node1441_r;
    reg node1441_l;
    reg node1442_r;
    reg node1442_l;
    reg node1443_r;
    reg node1443_l;
    reg node1444_r;
    reg node1444_l;
    reg node1445;
    reg node1446;
    reg node1447_r;
    reg node1447_l;
    reg node1448;
    reg node1449;
    reg node1450_r;
    reg node1450_l;
    reg node1451_r;
    reg node1451_l;
    reg node1452;
    reg node1453;
    reg node1454_r;
    reg node1454_l;
    reg node1455;
    reg node1456;
    reg node1457_r;
    reg node1457_l;
    reg node1458_r;
    reg node1458_l;
    reg node1459;
    reg node1460_r;
    reg node1460_l;
    reg node1461;
    reg node1462;
    reg node1463_r;
    reg node1463_l;
    reg node1464_r;
    reg node1464_l;
    reg node1465;
    reg node1466;
    reg node1467_r;
    reg node1467_l;
    reg node1468;
    reg node1469;
    reg node1470_r;
    reg node1470_l;
    reg node1471_r;
    reg node1471_l;
    reg node1472_r;
    reg node1472_l;
    reg node1473_r;
    reg node1473_l;
    reg node1474;
    reg node1475;
    reg node1476_r;
    reg node1476_l;
    reg node1477;
    reg node1478;
    reg node1479_r;
    reg node1479_l;
    reg node1480_r;
    reg node1480_l;
    reg node1481;
    reg node1482;
    reg node1483_r;
    reg node1483_l;
    reg node1484;
    reg node1485;
    reg node1486_r;
    reg node1486_l;
    reg node1487_r;
    reg node1487_l;
    reg node1488_r;
    reg node1488_l;
    reg node1489;
    reg node1490;
    reg node1491_r;
    reg node1491_l;
    reg node1492;
    reg node1493;
    reg node1494_r;
    reg node1494_l;
    reg node1495_r;
    reg node1495_l;
    reg node1496;
    reg node1497;
    reg node1498_r;
    reg node1498_l;
    reg node1499;
    reg node1500;
    reg node1501_r;
    reg node1501_l;
    reg node1502_r;
    reg node1502_l;
    reg node1503_r;
    reg node1503_l;
    reg node1504_r;
    reg node1504_l;
    reg node1505_r;
    reg node1505_l;
    reg node1506_r;
    reg node1506_l;
    reg node1507;
    reg node1508;
    reg node1509;
    reg node1510_r;
    reg node1510_l;
    reg node1511_r;
    reg node1511_l;
    reg node1512;
    reg node1513;
    reg node1514_r;
    reg node1514_l;
    reg node1515;
    reg node1516;
    reg node1517_r;
    reg node1517_l;
    reg node1518_r;
    reg node1518_l;
    reg node1519_r;
    reg node1519_l;
    reg node1520;
    reg node1521;
    reg node1522_r;
    reg node1522_l;
    reg node1523;
    reg node1524;
    reg node1525_r;
    reg node1525_l;
    reg node1526_r;
    reg node1526_l;
    reg node1527;
    reg node1528;
    reg node1529_r;
    reg node1529_l;
    reg node1530;
    reg node1531;
    reg node1532_r;
    reg node1532_l;
    reg node1533_r;
    reg node1533_l;
    reg node1534_r;
    reg node1534_l;
    reg node1535_r;
    reg node1535_l;
    reg node1536;
    reg node1537;
    reg node1538_r;
    reg node1538_l;
    reg node1539;
    reg node1540;
    reg node1541_r;
    reg node1541_l;
    reg node1542_r;
    reg node1542_l;
    reg node1543;
    reg node1544;
    reg node1545_r;
    reg node1545_l;
    reg node1546;
    reg node1547;
    reg node1548_r;
    reg node1548_l;
    reg node1549_r;
    reg node1549_l;
    reg node1550_r;
    reg node1550_l;
    reg node1551;
    reg node1552;
    reg node1553_r;
    reg node1553_l;
    reg node1554;
    reg node1555;
    reg node1556_r;
    reg node1556_l;
    reg node1557_r;
    reg node1557_l;
    reg node1558;
    reg node1559;
    reg node1560_r;
    reg node1560_l;
    reg node1561;
    reg node1562;
    reg node1563_r;
    reg node1563_l;
    reg node1564_r;
    reg node1564_l;
    reg node1565_r;
    reg node1565_l;
    reg node1566_r;
    reg node1566_l;
    reg node1567_r;
    reg node1567_l;
    reg node1568;
    reg node1569;
    reg node1570_r;
    reg node1570_l;
    reg node1571;
    reg node1572;
    reg node1573_r;
    reg node1573_l;
    reg node1574_r;
    reg node1574_l;
    reg node1575;
    reg node1576;
    reg node1577_r;
    reg node1577_l;
    reg node1578;
    reg node1579;
    reg node1580_r;
    reg node1580_l;
    reg node1581_r;
    reg node1581_l;
    reg node1582_r;
    reg node1582_l;
    reg node1583;
    reg node1584;
    reg node1585_r;
    reg node1585_l;
    reg node1586;
    reg node1587;
    reg node1588_r;
    reg node1588_l;
    reg node1589_r;
    reg node1589_l;
    reg node1590;
    reg node1591;
    reg node1592;
    reg node1593_r;
    reg node1593_l;
    reg node1594_r;
    reg node1594_l;
    reg node1595_r;
    reg node1595_l;
    reg node1596_r;
    reg node1596_l;
    reg node1597;
    reg node1598;
    reg node1599_r;
    reg node1599_l;
    reg node1600;
    reg node1601;
    reg node1602_r;
    reg node1602_l;
    reg node1603_r;
    reg node1603_l;
    reg node1604;
    reg node1605;
    reg node1606_r;
    reg node1606_l;
    reg node1607;
    reg node1608;
    reg node1609_r;
    reg node1609_l;
    reg node1610_r;
    reg node1610_l;
    reg node1611_r;
    reg node1611_l;
    reg node1612;
    reg node1613;
    reg node1614_r;
    reg node1614_l;
    reg node1615;
    reg node1616;
    reg node1617_r;
    reg node1617_l;
    reg node1618_r;
    reg node1618_l;
    reg node1619;
    reg node1620;
    reg node1621_r;
    reg node1621_l;
    reg node1622;
    reg node1623;
    reg node1624_r;
    reg node1624_l;
    reg node1625_r;
    reg node1625_l;
    reg node1626_r;
    reg node1626_l;
    reg node1627_r;
    reg node1627_l;
    reg node1628_r;
    reg node1628_l;
    reg node1629_r;
    reg node1629_l;
    reg node1630_r;
    reg node1630_l;
    reg node1631;
    reg node1632;
    reg node1633;
    reg node1634_r;
    reg node1634_l;
    reg node1635_r;
    reg node1635_l;
    reg node1636;
    reg node1637;
    reg node1638_r;
    reg node1638_l;
    reg node1639;
    reg node1640;
    reg node1641_r;
    reg node1641_l;
    reg node1642_r;
    reg node1642_l;
    reg node1643_r;
    reg node1643_l;
    reg node1644;
    reg node1645;
    reg node1646_r;
    reg node1646_l;
    reg node1647;
    reg node1648;
    reg node1649_r;
    reg node1649_l;
    reg node1650;
    reg node1651_r;
    reg node1651_l;
    reg node1652;
    reg node1653;
    reg node1654_r;
    reg node1654_l;
    reg node1655_r;
    reg node1655_l;
    reg node1656_r;
    reg node1656_l;
    reg node1657_r;
    reg node1657_l;
    reg node1658;
    reg node1659;
    reg node1660_r;
    reg node1660_l;
    reg node1661;
    reg node1662;
    reg node1663_r;
    reg node1663_l;
    reg node1664_r;
    reg node1664_l;
    reg node1665;
    reg node1666;
    reg node1667_r;
    reg node1667_l;
    reg node1668;
    reg node1669;
    reg node1670_r;
    reg node1670_l;
    reg node1671_r;
    reg node1671_l;
    reg node1672_r;
    reg node1672_l;
    reg node1673;
    reg node1674;
    reg node1675_r;
    reg node1675_l;
    reg node1676;
    reg node1677;
    reg node1678_r;
    reg node1678_l;
    reg node1679;
    reg node1680;
    reg node1681_r;
    reg node1681_l;
    reg node1682_r;
    reg node1682_l;
    reg node1683_r;
    reg node1683_l;
    reg node1684_r;
    reg node1684_l;
    reg node1685_r;
    reg node1685_l;
    reg node1686;
    reg node1687;
    reg node1688_r;
    reg node1688_l;
    reg node1689;
    reg node1690;
    reg node1691_r;
    reg node1691_l;
    reg node1692_r;
    reg node1692_l;
    reg node1693;
    reg node1694;
    reg node1695;
    reg node1696_r;
    reg node1696_l;
    reg node1697_r;
    reg node1697_l;
    reg node1698_r;
    reg node1698_l;
    reg node1699;
    reg node1700;
    reg node1701_r;
    reg node1701_l;
    reg node1702;
    reg node1703;
    reg node1704_r;
    reg node1704_l;
    reg node1705_r;
    reg node1705_l;
    reg node1706;
    reg node1707;
    reg node1708_r;
    reg node1708_l;
    reg node1709;
    reg node1710;
    reg node1711_r;
    reg node1711_l;
    reg node1712_r;
    reg node1712_l;
    reg node1713_r;
    reg node1713_l;
    reg node1714_r;
    reg node1714_l;
    reg node1715;
    reg node1716;
    reg node1717_r;
    reg node1717_l;
    reg node1718;
    reg node1719;
    reg node1720_r;
    reg node1720_l;
    reg node1721_r;
    reg node1721_l;
    reg node1722;
    reg node1723;
    reg node1724_r;
    reg node1724_l;
    reg node1725;
    reg node1726;
    reg node1727_r;
    reg node1727_l;
    reg node1728_r;
    reg node1728_l;
    reg node1729;
    reg node1730_r;
    reg node1730_l;
    reg node1731;
    reg node1732;
    reg node1733_r;
    reg node1733_l;
    reg node1734_r;
    reg node1734_l;
    reg node1735;
    reg node1736;
    reg node1737_r;
    reg node1737_l;
    reg node1738;
    reg node1739;
    reg node1740_r;
    reg node1740_l;
    reg node1741_r;
    reg node1741_l;
    reg node1742_r;
    reg node1742_l;
    reg node1743_r;
    reg node1743_l;
    reg node1744_r;
    reg node1744_l;
    reg node1745_r;
    reg node1745_l;
    reg node1746;
    reg node1747;
    reg node1748_r;
    reg node1748_l;
    reg node1749;
    reg node1750;
    reg node1751_r;
    reg node1751_l;
    reg node1752_r;
    reg node1752_l;
    reg node1753;
    reg node1754;
    reg node1755_r;
    reg node1755_l;
    reg node1756;
    reg node1757;
    reg node1758_r;
    reg node1758_l;
    reg node1759_r;
    reg node1759_l;
    reg node1760;
    reg node1761;
    reg node1762_r;
    reg node1762_l;
    reg node1763;
    reg node1764;
    reg node1765_r;
    reg node1765_l;
    reg node1766_r;
    reg node1766_l;
    reg node1767_r;
    reg node1767_l;
    reg node1768_r;
    reg node1768_l;
    reg node1769;
    reg node1770;
    reg node1771_r;
    reg node1771_l;
    reg node1772;
    reg node1773;
    reg node1774_r;
    reg node1774_l;
    reg node1775_r;
    reg node1775_l;
    reg node1776;
    reg node1777;
    reg node1778;
    reg node1779_r;
    reg node1779_l;
    reg node1780;
    reg node1781;
    reg node1782_r;
    reg node1782_l;
    reg node1783_r;
    reg node1783_l;
    reg node1784_r;
    reg node1784_l;
    reg node1785;
    reg node1786_r;
    reg node1786_l;
    reg node1787;
    reg node1788;
    reg node1789_r;
    reg node1789_l;
    reg node1790_r;
    reg node1790_l;
    reg node1791_r;
    reg node1791_l;
    reg node1792;
    reg node1793;
    reg node1794_r;
    reg node1794_l;
    reg node1795;
    reg node1796;
    reg node1797_r;
    reg node1797_l;
    reg node1798_r;
    reg node1798_l;
    reg node1799;
    reg node1800;
    reg node1801_r;
    reg node1801_l;
    reg node1802;
    reg node1803;
    reg node1804_r;
    reg node1804_l;
    reg node1805_r;
    reg node1805_l;
    reg node1806_r;
    reg node1806_l;
    reg node1807_r;
    reg node1807_l;
    reg node1808;
    reg node1809;
    reg node1810_r;
    reg node1810_l;
    reg node1811;
    reg node1812;
    reg node1813_r;
    reg node1813_l;
    reg node1814_r;
    reg node1814_l;
    reg node1815;
    reg node1816;
    reg node1817_r;
    reg node1817_l;
    reg node1818;
    reg node1819;
    reg node1820_r;
    reg node1820_l;
    reg node1821_r;
    reg node1821_l;
    reg node1822;
    reg node1823_r;
    reg node1823_l;
    reg node1824;
    reg node1825;
    reg node1826_r;
    reg node1826_l;
    reg node1827_r;
    reg node1827_l;
    reg node1828;
    reg node1829;
    reg node1830;
    reg result0;
    reg result1;
    reg result2;
    reg result3;
    reg result4;
    reg result5;
    reg result6;
    reg result7;
    reg result8;
    reg result9;

    begin
      node0_r = pixel[155];
      node0_l = ~pixel[155];
      node1_r = node0_l & pixel[263];
      node1_l = node0_l & ~pixel[263];
      node2_r = node1_l & pixel[322];
      node2_l = node1_l & ~pixel[322];
      node3_r = node2_l & pixel[400];
      node3_l = node2_l & ~pixel[400];
      node4_r = node3_l & pixel[239];
      node4_l = node3_l & ~pixel[239];
      node5_r = node4_l & pixel[624];
      node5_l = node4_l & ~pixel[624];
      node6_r = node5_l & pixel[571];
      node6_l = node5_l & ~pixel[571];
      node7_r = node6_l & pixel[209];
      node7_l = node6_l & ~pixel[209];
      node8_r = node7_l & pixel[350];
      node8_l = node7_l & ~pixel[350];
      node9_r = node8_l & pixel[524];
      node9_l = node8_l & ~pixel[524];
      node10 = node9_l;
      node11 = node9_r;
      node12_r = node8_r & pixel[205];
      node12_l = node8_r & ~pixel[205];
      node13 = node12_l;
      node14 = node12_r;
      node15_r = node7_r & pixel[426];
      node15_l = node7_r & ~pixel[426];
      node16_r = node15_l & pixel[320];
      node16_l = node15_l & ~pixel[320];
      node17 = node16_l;
      node18 = node16_r;
      node19_r = node15_r & pixel[569];
      node19_l = node15_r & ~pixel[569];
      node20 = node19_l;
      node21 = node19_r;
      node22_r = node6_r & pixel[269];
      node22_l = node6_r & ~pixel[269];
      node23_r = node22_l & pixel[369];
      node23_l = node22_l & ~pixel[369];
      node24_r = node23_l & pixel[601];
      node24_l = node23_l & ~pixel[601];
      node25 = node24_l;
      node26 = node24_r;
      node27_r = node23_r & pixel[632];
      node27_l = node23_r & ~pixel[632];
      node28 = node27_l;
      node29 = node27_r;
      node30_r = node22_r & pixel[433];
      node30_l = node22_r & ~pixel[433];
      node31_r = node30_l & pixel[219];
      node31_l = node30_l & ~pixel[219];
      node32 = node31_l;
      node33 = node31_r;
      node34_r = node30_r & pixel[374];
      node34_l = node30_r & ~pixel[374];
      node35 = node34_l;
      node36 = node34_r;
      node37_r = node5_r & pixel[101];
      node37_l = node5_r & ~pixel[101];
      node38_r = node37_l & pixel[488];
      node38_l = node37_l & ~pixel[488];
      node39_r = node38_l & pixel[265];
      node39_l = node38_l & ~pixel[265];
      node40_r = node39_l & pixel[471];
      node40_l = node39_l & ~pixel[471];
      node41 = node40_l;
      node42 = node40_r;
      node43_r = node39_r & pixel[482];
      node43_l = node39_r & ~pixel[482];
      node44 = node43_l;
      node45 = node43_r;
      node46_r = node38_r & pixel[234];
      node46_l = node38_r & ~pixel[234];
      node47_r = node46_l & pixel[430];
      node47_l = node46_l & ~pixel[430];
      node48 = node47_l;
      node49 = node47_r;
      node50_r = node46_r & pixel[629];
      node50_l = node46_r & ~pixel[629];
      node51 = node50_l;
      node52 = node50_r;
      node53_r = node37_r & pixel[323];
      node53_l = node37_r & ~pixel[323];
      node54_r = node53_l & pixel[228];
      node54_l = node53_l & ~pixel[228];
      node55_r = node54_l & pixel[347];
      node55_l = node54_l & ~pixel[347];
      node56 = node55_l;
      node57 = node55_r;
      node58 = node54_r;
      node59_r = node53_r & pixel[461];
      node59_l = node53_r & ~pixel[461];
      node60 = node59_l;
      node61_r = node59_r & pixel[628];
      node61_l = node59_r & ~pixel[628];
      node62 = node61_l;
      node63 = node61_r;
      node64_r = node4_r & pixel[291];
      node64_l = node4_r & ~pixel[291];
      node65_r = node64_l & pixel[433];
      node65_l = node64_l & ~pixel[433];
      node66_r = node65_l & pixel[208];
      node66_l = node65_l & ~pixel[208];
      node67_r = node66_l & pixel[192];
      node67_l = node66_l & ~pixel[192];
      node68_r = node67_l & pixel[416];
      node68_l = node67_l & ~pixel[416];
      node69 = node68_l;
      node70 = node68_r;
      node71 = node67_r;
      node72_r = node66_r & pixel[454];
      node72_l = node66_r & ~pixel[454];
      node73_r = node72_l & pixel[577];
      node73_l = node72_l & ~pixel[577];
      node74 = node73_l;
      node75 = node73_r;
      node76_r = node72_r & pixel[600];
      node76_l = node72_r & ~pixel[600];
      node77 = node76_l;
      node78 = node76_r;
      node79_r = node65_r & pixel[544];
      node79_l = node65_r & ~pixel[544];
      node80_r = node79_l & pixel[209];
      node80_l = node79_l & ~pixel[209];
      node81_r = node80_l & pixel[553];
      node81_l = node80_l & ~pixel[553];
      node82 = node81_l;
      node83 = node81_r;
      node84_r = node80_r & pixel[488];
      node84_l = node80_r & ~pixel[488];
      node85 = node84_l;
      node86 = node84_r;
      node87_r = node79_r & pixel[344];
      node87_l = node79_r & ~pixel[344];
      node88_r = node87_l & pixel[709];
      node88_l = node87_l & ~pixel[709];
      node89 = node88_l;
      node90 = node88_r;
      node91 = node87_r;
      node92_r = node64_r & pixel[566];
      node92_l = node64_r & ~pixel[566];
      node93_r = node92_l & pixel[569];
      node93_l = node92_l & ~pixel[569];
      node94_r = node93_l & pixel[623];
      node94_l = node93_l & ~pixel[623];
      node95_r = node94_l & pixel[343];
      node95_l = node94_l & ~pixel[343];
      node96 = node95_l;
      node97 = node95_r;
      node98 = node94_r;
      node99_r = node93_r & pixel[103];
      node99_l = node93_r & ~pixel[103];
      node100_r = node99_l & pixel[354];
      node100_l = node99_l & ~pixel[354];
      node101 = node100_l;
      node102 = node100_r;
      node103_r = node99_r & pixel[430];
      node103_l = node99_r & ~pixel[430];
      node104 = node103_l;
      node105 = node103_r;
      node106_r = node92_r & pixel[513];
      node106_l = node92_r & ~pixel[513];
      node107_r = node106_l & pixel[412];
      node107_l = node106_l & ~pixel[412];
      node108_r = node107_l & pixel[356];
      node108_l = node107_l & ~pixel[356];
      node109 = node108_l;
      node110 = node108_r;
      node111_r = node107_r & pixel[133];
      node111_l = node107_r & ~pixel[133];
      node112 = node111_l;
      node113 = node111_r;
      node114_r = node106_r & pixel[624];
      node114_l = node106_r & ~pixel[624];
      node115_r = node114_l & pixel[535];
      node115_l = node114_l & ~pixel[535];
      node116 = node115_l;
      node117 = node115_r;
      node118 = node114_r;
      node119_r = node3_r & pixel[571];
      node119_l = node3_r & ~pixel[571];
      node120_r = node119_l & pixel[653];
      node120_l = node119_l & ~pixel[653];
      node121_r = node120_l & pixel[240];
      node121_l = node120_l & ~pixel[240];
      node122_r = node121_l & pixel[96];
      node122_l = node121_l & ~pixel[96];
      node123_r = node122_l & pixel[65];
      node123_l = node122_l & ~pixel[65];
      node124_r = node123_l & pixel[216];
      node124_l = node123_l & ~pixel[216];
      node125 = node124_l;
      node126 = node124_r;
      node127 = node123_r;
      node128_r = node122_r & pixel[302];
      node128_l = node122_r & ~pixel[302];
      node129 = node128_l;
      node130_r = node128_r & pixel[381];
      node130_l = node128_r & ~pixel[381];
      node131 = node130_l;
      node132 = node130_r;
      node133_r = node121_r & pixel[181];
      node133_l = node121_r & ~pixel[181];
      node134_r = node133_l & pixel[239];
      node134_l = node133_l & ~pixel[239];
      node135_r = node134_l & pixel[190];
      node135_l = node134_l & ~pixel[190];
      node136 = node135_l;
      node137 = node135_r;
      node138_r = node134_r & pixel[373];
      node138_l = node134_r & ~pixel[373];
      node139 = node138_l;
      node140 = node138_r;
      node141_r = node133_r & pixel[521];
      node141_l = node133_r & ~pixel[521];
      node142_r = node141_l & pixel[569];
      node142_l = node141_l & ~pixel[569];
      node143 = node142_l;
      node144 = node142_r;
      node145_r = node141_r & pixel[287];
      node145_l = node141_r & ~pixel[287];
      node146 = node145_l;
      node147 = node145_r;
      node148_r = node120_r & pixel[509];
      node148_l = node120_r & ~pixel[509];
      node149_r = node148_l & pixel[298];
      node149_l = node148_l & ~pixel[298];
      node150_r = node149_l & pixel[191];
      node150_l = node149_l & ~pixel[191];
      node151_r = node150_l & pixel[511];
      node151_l = node150_l & ~pixel[511];
      node152 = node151_l;
      node153 = node151_r;
      node154 = node150_r;
      node155_r = node149_r & pixel[374];
      node155_l = node149_r & ~pixel[374];
      node156_r = node155_l & pixel[380];
      node156_l = node155_l & ~pixel[380];
      node157 = node156_l;
      node158 = node156_r;
      node159_r = node155_r & pixel[711];
      node159_l = node155_r & ~pixel[711];
      node160 = node159_l;
      node161 = node159_r;
      node162_r = node148_r & pixel[539];
      node162_l = node148_r & ~pixel[539];
      node163_r = node162_l & pixel[214];
      node163_l = node162_l & ~pixel[214];
      node164 = node163_l;
      node165_r = node163_r & pixel[660];
      node165_l = node163_r & ~pixel[660];
      node166 = node165_l;
      node167 = node165_r;
      node168 = node162_r;
      node169_r = node119_r & pixel[123];
      node169_l = node119_r & ~pixel[123];
      node170_r = node169_l & pixel[120];
      node170_l = node169_l & ~pixel[120];
      node171_r = node170_l & pixel[538];
      node171_l = node170_l & ~pixel[538];
      node172_r = node171_l & pixel[238];
      node172_l = node171_l & ~pixel[238];
      node173_r = node172_l & pixel[71];
      node173_l = node172_l & ~pixel[71];
      node174 = node173_l;
      node175 = node173_r;
      node176_r = node172_r & pixel[381];
      node176_l = node172_r & ~pixel[381];
      node177 = node176_l;
      node178 = node176_r;
      node179_r = node171_r & pixel[377];
      node179_l = node171_r & ~pixel[377];
      node180_r = node179_l & pixel[626];
      node180_l = node179_l & ~pixel[626];
      node181 = node180_l;
      node182 = node180_r;
      node183_r = node179_r & pixel[320];
      node183_l = node179_r & ~pixel[320];
      node184 = node183_l;
      node185 = node183_r;
      node186_r = node170_r & pixel[153];
      node186_l = node170_r & ~pixel[153];
      node187_r = node186_l & pixel[214];
      node187_l = node186_l & ~pixel[214];
      node188_r = node187_l & pixel[574];
      node188_l = node187_l & ~pixel[574];
      node189 = node188_l;
      node190 = node188_r;
      node191 = node187_r;
      node192 = node186_r;
      node193_r = node169_r & pixel[268];
      node193_l = node169_r & ~pixel[268];
      node194_r = node193_l & pixel[130];
      node194_l = node193_l & ~pixel[130];
      node195_r = node194_l & pixel[245];
      node195_l = node194_l & ~pixel[245];
      node196_r = node195_l & pixel[403];
      node196_l = node195_l & ~pixel[403];
      node197 = node196_l;
      node198 = node196_r;
      node199_r = node195_r & pixel[407];
      node199_l = node195_r & ~pixel[407];
      node200 = node199_l;
      node201 = node199_r;
      node202_r = node194_r & pixel[344];
      node202_l = node194_r & ~pixel[344];
      node203 = node202_l;
      node204_r = node202_r & pixel[300];
      node204_l = node202_r & ~pixel[300];
      node205 = node204_l;
      node206 = node204_r;
      node207_r = node193_r & pixel[521];
      node207_l = node193_r & ~pixel[521];
      node208_r = node207_l & pixel[404];
      node208_l = node207_l & ~pixel[404];
      node209_r = node208_l & pixel[260];
      node209_l = node208_l & ~pixel[260];
      node210 = node209_l;
      node211 = node209_r;
      node212_r = node208_r & pixel[413];
      node212_l = node208_r & ~pixel[413];
      node213 = node212_l;
      node214 = node212_r;
      node215_r = node207_r & pixel[237];
      node215_l = node207_r & ~pixel[237];
      node216 = node215_l;
      node217 = node215_r;
      node218_r = node2_r & pixel[430];
      node218_l = node2_r & ~pixel[430];
      node219_r = node218_l & pixel[347];
      node219_l = node218_l & ~pixel[347];
      node220_r = node219_l & pixel[550];
      node220_l = node219_l & ~pixel[550];
      node221_r = node220_l & pixel[466];
      node221_l = node220_l & ~pixel[466];
      node222_r = node221_l & pixel[204];
      node222_l = node221_l & ~pixel[204];
      node223_r = node222_l & pixel[454];
      node223_l = node222_l & ~pixel[454];
      node224_r = node223_l & pixel[409];
      node224_l = node223_l & ~pixel[409];
      node225 = node224_l;
      node226 = node224_r;
      node227_r = node223_r & pixel[541];
      node227_l = node223_r & ~pixel[541];
      node228 = node227_l;
      node229 = node227_r;
      node230_r = node222_r & pixel[607];
      node230_l = node222_r & ~pixel[607];
      node231_r = node230_l & pixel[380];
      node231_l = node230_l & ~pixel[380];
      node232 = node231_l;
      node233 = node231_r;
      node234_r = node230_r & pixel[358];
      node234_l = node230_r & ~pixel[358];
      node235 = node234_l;
      node236 = node234_r;
      node237_r = node221_r & pixel[486];
      node237_l = node221_r & ~pixel[486];
      node238_r = node237_l & pixel[291];
      node238_l = node237_l & ~pixel[291];
      node239_r = node238_l & pixel[461];
      node239_l = node238_l & ~pixel[461];
      node240 = node239_l;
      node241 = node239_r;
      node242_r = node238_r & pixel[384];
      node242_l = node238_r & ~pixel[384];
      node243 = node242_l;
      node244 = node242_r;
      node245_r = node237_r & pixel[710];
      node245_l = node237_r & ~pixel[710];
      node246_r = node245_l & pixel[102];
      node246_l = node245_l & ~pixel[102];
      node247 = node246_l;
      node248 = node246_r;
      node249 = node245_r;
      node250_r = node220_r & pixel[370];
      node250_l = node220_r & ~pixel[370];
      node251_r = node250_l & pixel[518];
      node251_l = node250_l & ~pixel[518];
      node252_r = node251_l & pixel[319];
      node252_l = node251_l & ~pixel[319];
      node253_r = node252_l & pixel[517];
      node253_l = node252_l & ~pixel[517];
      node254 = node253_l;
      node255 = node253_r;
      node256_r = node252_r & pixel[352];
      node256_l = node252_r & ~pixel[352];
      node257 = node256_l;
      node258 = node256_r;
      node259_r = node251_r & pixel[414];
      node259_l = node251_r & ~pixel[414];
      node260_r = node259_l & pixel[152];
      node260_l = node259_l & ~pixel[152];
      node261 = node260_l;
      node262 = node260_r;
      node263_r = node259_r & pixel[471];
      node263_l = node259_r & ~pixel[471];
      node264 = node263_l;
      node265 = node263_r;
      node266_r = node250_r & pixel[405];
      node266_l = node250_r & ~pixel[405];
      node267_r = node266_l & pixel[512];
      node267_l = node266_l & ~pixel[512];
      node268_r = node267_l & pixel[240];
      node268_l = node267_l & ~pixel[240];
      node269 = node268_l;
      node270 = node268_r;
      node271_r = node267_r & pixel[344];
      node271_l = node267_r & ~pixel[344];
      node272 = node271_l;
      node273 = node271_r;
      node274_r = node266_r & pixel[189];
      node274_l = node266_r & ~pixel[189];
      node275_r = node274_l & pixel[574];
      node275_l = node274_l & ~pixel[574];
      node276 = node275_l;
      node277 = node275_r;
      node278 = node274_r;
      node279_r = node219_r & pixel[210];
      node279_l = node219_r & ~pixel[210];
      node280_r = node279_l & pixel[539];
      node280_l = node279_l & ~pixel[539];
      node281_r = node280_l & pixel[177];
      node281_l = node280_l & ~pixel[177];
      node282_r = node281_l & pixel[565];
      node282_l = node281_l & ~pixel[565];
      node283_r = node282_l & pixel[318];
      node283_l = node282_l & ~pixel[318];
      node284 = node283_l;
      node285 = node283_r;
      node286_r = node282_r & pixel[413];
      node286_l = node282_r & ~pixel[413];
      node287 = node286_l;
      node288 = node286_r;
      node289_r = node281_r & pixel[497];
      node289_l = node281_r & ~pixel[497];
      node290_r = node289_l & pixel[607];
      node290_l = node289_l & ~pixel[607];
      node291 = node290_l;
      node292 = node290_r;
      node293_r = node289_r & pixel[243];
      node293_l = node289_r & ~pixel[243];
      node294 = node293_l;
      node295 = node293_r;
      node296_r = node280_r & pixel[469];
      node296_l = node280_r & ~pixel[469];
      node297_r = node296_l & pixel[441];
      node297_l = node296_l & ~pixel[441];
      node298_r = node297_l & pixel[467];
      node298_l = node297_l & ~pixel[467];
      node299 = node298_l;
      node300 = node298_r;
      node301_r = node297_r & pixel[244];
      node301_l = node297_r & ~pixel[244];
      node302 = node301_l;
      node303 = node301_r;
      node304_r = node296_r & pixel[414];
      node304_l = node296_r & ~pixel[414];
      node305 = node304_l;
      node306_r = node304_r & pixel[461];
      node306_l = node304_r & ~pixel[461];
      node307 = node306_l;
      node308 = node306_r;
      node309_r = node279_r & pixel[219];
      node309_l = node279_r & ~pixel[219];
      node310_r = node309_l & pixel[260];
      node310_l = node309_l & ~pixel[260];
      node311_r = node310_l & pixel[573];
      node311_l = node310_l & ~pixel[573];
      node312_r = node311_l & pixel[185];
      node312_l = node311_l & ~pixel[185];
      node313 = node312_l;
      node314 = node312_r;
      node315_r = node311_r & pixel[204];
      node315_l = node311_r & ~pixel[204];
      node316 = node315_l;
      node317 = node315_r;
      node318_r = node310_r & pixel[492];
      node318_l = node310_r & ~pixel[492];
      node319_r = node318_l & pixel[287];
      node319_l = node318_l & ~pixel[287];
      node320 = node319_l;
      node321 = node319_r;
      node322_r = node318_r & pixel[203];
      node322_l = node318_r & ~pixel[203];
      node323 = node322_l;
      node324 = node322_r;
      node325_r = node309_r & pixel[329];
      node325_l = node309_r & ~pixel[329];
      node326_r = node325_l & pixel[216];
      node326_l = node325_l & ~pixel[216];
      node327_r = node326_l & pixel[594];
      node327_l = node326_l & ~pixel[594];
      node328 = node327_l;
      node329 = node327_r;
      node330_r = node326_r & pixel[202];
      node330_l = node326_r & ~pixel[202];
      node331 = node330_l;
      node332 = node330_r;
      node333_r = node325_r & pixel[386];
      node333_l = node325_r & ~pixel[386];
      node334_r = node333_l & pixel[511];
      node334_l = node333_l & ~pixel[511];
      node335 = node334_l;
      node336 = node334_r;
      node337_r = node333_r & pixel[399];
      node337_l = node333_r & ~pixel[399];
      node338 = node337_l;
      node339 = node337_r;
      node340_r = node218_r & pixel[594];
      node340_l = node218_r & ~pixel[594];
      node341_r = node340_l & pixel[186];
      node341_l = node340_l & ~pixel[186];
      node342_r = node341_l & pixel[524];
      node342_l = node341_l & ~pixel[524];
      node343_r = node342_l & pixel[181];
      node343_l = node342_l & ~pixel[181];
      node344_r = node343_l & pixel[410];
      node344_l = node343_l & ~pixel[410];
      node345_r = node344_l & pixel[296];
      node345_l = node344_l & ~pixel[296];
      node346 = node345_l;
      node347 = node345_r;
      node348_r = node344_r & pixel[539];
      node348_l = node344_r & ~pixel[539];
      node349 = node348_l;
      node350 = node348_r;
      node351_r = node343_r & pixel[314];
      node351_l = node343_r & ~pixel[314];
      node352_r = node351_l & pixel[122];
      node352_l = node351_l & ~pixel[122];
      node353 = node352_l;
      node354 = node352_r;
      node355_r = node351_r & pixel[233];
      node355_l = node351_r & ~pixel[233];
      node356 = node355_l;
      node357 = node355_r;
      node358_r = node342_r & pixel[572];
      node358_l = node342_r & ~pixel[572];
      node359_r = node358_l & pixel[178];
      node359_l = node358_l & ~pixel[178];
      node360_r = node359_l & pixel[271];
      node360_l = node359_l & ~pixel[271];
      node361 = node360_l;
      node362 = node360_r;
      node363_r = node359_r & pixel[519];
      node363_l = node359_r & ~pixel[519];
      node364 = node363_l;
      node365 = node363_r;
      node366_r = node358_r & pixel[386];
      node366_l = node358_r & ~pixel[386];
      node367_r = node366_l & pixel[660];
      node367_l = node366_l & ~pixel[660];
      node368 = node367_l;
      node369 = node367_r;
      node370_r = node366_r & pixel[238];
      node370_l = node366_r & ~pixel[238];
      node371 = node370_l;
      node372 = node370_r;
      node373_r = node341_r & pixel[105];
      node373_l = node341_r & ~pixel[105];
      node374_r = node373_l & pixel[101];
      node374_l = node373_l & ~pixel[101];
      node375_r = node374_l & pixel[353];
      node375_l = node374_l & ~pixel[353];
      node376_r = node375_l & pixel[328];
      node376_l = node375_l & ~pixel[328];
      node377 = node376_l;
      node378 = node376_r;
      node379_r = node375_r & pixel[347];
      node379_l = node375_r & ~pixel[347];
      node380 = node379_l;
      node381 = node379_r;
      node382_r = node374_r & pixel[99];
      node382_l = node374_r & ~pixel[99];
      node383_r = node382_l & pixel[156];
      node383_l = node382_l & ~pixel[156];
      node384 = node383_l;
      node385 = node383_r;
      node386_r = node382_r & pixel[265];
      node386_l = node382_r & ~pixel[265];
      node387 = node386_l;
      node388 = node386_r;
      node389_r = node373_r & pixel[425];
      node389_l = node373_r & ~pixel[425];
      node390_r = node389_l & pixel[597];
      node390_l = node389_l & ~pixel[597];
      node391_r = node390_l & pixel[549];
      node391_l = node390_l & ~pixel[549];
      node392 = node391_l;
      node393 = node391_r;
      node394_r = node390_r & pixel[439];
      node394_l = node390_r & ~pixel[439];
      node395 = node394_l;
      node396 = node394_r;
      node397 = node389_r;
      node398_r = node340_r & pixel[384];
      node398_l = node340_r & ~pixel[384];
      node399_r = node398_l & pixel[213];
      node399_l = node398_l & ~pixel[213];
      node400_r = node399_l & pixel[649];
      node400_l = node399_l & ~pixel[649];
      node401_r = node400_l & pixel[133];
      node401_l = node400_l & ~pixel[133];
      node402_r = node401_l & pixel[497];
      node402_l = node401_l & ~pixel[497];
      node403 = node402_l;
      node404 = node402_r;
      node405_r = node401_r & pixel[437];
      node405_l = node401_r & ~pixel[437];
      node406 = node405_l;
      node407 = node405_r;
      node408_r = node400_r & pixel[573];
      node408_l = node400_r & ~pixel[573];
      node409 = node408_l;
      node410 = node408_r;
      node411_r = node399_r & pixel[386];
      node411_l = node399_r & ~pixel[386];
      node412_r = node411_l & pixel[328];
      node412_l = node411_l & ~pixel[328];
      node413_r = node412_l & pixel[347];
      node413_l = node412_l & ~pixel[347];
      node414 = node413_l;
      node415 = node413_r;
      node416_r = node412_r & pixel[296];
      node416_l = node412_r & ~pixel[296];
      node417 = node416_l;
      node418 = node416_r;
      node419 = node411_r;
      node420_r = node398_r & pixel[467];
      node420_l = node398_r & ~pixel[467];
      node421_r = node420_l & pixel[458];
      node421_l = node420_l & ~pixel[458];
      node422_r = node421_l & pixel[235];
      node422_l = node421_l & ~pixel[235];
      node423_r = node422_l & pixel[301];
      node423_l = node422_l & ~pixel[301];
      node424 = node423_l;
      node425 = node423_r;
      node426 = node422_r;
      node427_r = node421_r & pixel[460];
      node427_l = node421_r & ~pixel[460];
      node428_r = node427_l & pixel[493];
      node428_l = node427_l & ~pixel[493];
      node429 = node428_l;
      node430 = node428_r;
      node431_r = node427_r & pixel[489];
      node431_l = node427_r & ~pixel[489];
      node432 = node431_l;
      node433 = node431_r;
      node434_r = node420_r & pixel[488];
      node434_l = node420_r & ~pixel[488];
      node435_r = node434_l & pixel[207];
      node435_l = node434_l & ~pixel[207];
      node436_r = node435_l & pixel[105];
      node436_l = node435_l & ~pixel[105];
      node437 = node436_l;
      node438 = node436_r;
      node439 = node435_r;
      node440_r = node434_r & pixel[246];
      node440_l = node434_r & ~pixel[246];
      node441_r = node440_l & pixel[607];
      node441_l = node440_l & ~pixel[607];
      node442 = node441_l;
      node443 = node441_r;
      node444_r = node440_r & pixel[348];
      node444_l = node440_r & ~pixel[348];
      node445 = node444_l;
      node446 = node444_r;
      node447_r = node1_r & pixel[429];
      node447_l = node1_r & ~pixel[429];
      node448_r = node447_l & pixel[405];
      node448_l = node447_l & ~pixel[405];
      node449_r = node448_l & pixel[387];
      node449_l = node448_l & ~pixel[387];
      node450_r = node449_l & pixel[566];
      node450_l = node449_l & ~pixel[566];
      node451_r = node450_l & pixel[553];
      node451_l = node450_l & ~pixel[553];
      node452_r = node451_l & pixel[454];
      node452_l = node451_l & ~pixel[454];
      node453_r = node452_l & pixel[374];
      node453_l = node452_l & ~pixel[374];
      node454_r = node453_l & pixel[150];
      node454_l = node453_l & ~pixel[150];
      node455 = node454_l;
      node456 = node454_r;
      node457_r = node453_r & pixel[294];
      node457_l = node453_r & ~pixel[294];
      node458 = node457_l;
      node459 = node457_r;
      node460_r = node452_r & pixel[516];
      node460_l = node452_r & ~pixel[516];
      node461_r = node460_l & pixel[489];
      node461_l = node460_l & ~pixel[489];
      node462 = node461_l;
      node463 = node461_r;
      node464_r = node460_r & pixel[210];
      node464_l = node460_r & ~pixel[210];
      node465 = node464_l;
      node466 = node464_r;
      node467_r = node451_r & pixel[555];
      node467_l = node451_r & ~pixel[555];
      node468_r = node467_l & pixel[257];
      node468_l = node467_l & ~pixel[257];
      node469_r = node468_l & pixel[454];
      node469_l = node468_l & ~pixel[454];
      node470 = node469_l;
      node471 = node469_r;
      node472_r = node468_r & pixel[178];
      node472_l = node468_r & ~pixel[178];
      node473 = node472_l;
      node474 = node472_r;
      node475_r = node467_r & pixel[441];
      node475_l = node467_r & ~pixel[441];
      node476_r = node475_l & pixel[691];
      node476_l = node475_l & ~pixel[691];
      node477 = node476_l;
      node478 = node476_r;
      node479_r = node475_r & pixel[236];
      node479_l = node475_r & ~pixel[236];
      node480 = node479_l;
      node481 = node479_r;
      node482_r = node450_r & pixel[349];
      node482_l = node450_r & ~pixel[349];
      node483_r = node482_l & pixel[629];
      node483_l = node482_l & ~pixel[629];
      node484_r = node483_l & pixel[655];
      node484_l = node483_l & ~pixel[655];
      node485_r = node484_l & pixel[134];
      node485_l = node484_l & ~pixel[134];
      node486 = node485_l;
      node487 = node485_r;
      node488_r = node484_r & pixel[513];
      node488_l = node484_r & ~pixel[513];
      node489 = node488_l;
      node490 = node488_r;
      node491_r = node483_r & pixel[496];
      node491_l = node483_r & ~pixel[496];
      node492_r = node491_l & pixel[328];
      node492_l = node491_l & ~pixel[328];
      node493 = node492_l;
      node494 = node492_r;
      node495_r = node491_r & pixel[485];
      node495_l = node491_r & ~pixel[485];
      node496 = node495_l;
      node497 = node495_r;
      node498_r = node482_r & pixel[620];
      node498_l = node482_r & ~pixel[620];
      node499_r = node498_l & pixel[414];
      node499_l = node498_l & ~pixel[414];
      node500_r = node499_l & pixel[380];
      node500_l = node499_l & ~pixel[380];
      node501 = node500_l;
      node502 = node500_r;
      node503_r = node499_r & pixel[683];
      node503_l = node499_r & ~pixel[683];
      node504 = node503_l;
      node505 = node503_r;
      node506_r = node498_r & pixel[709];
      node506_l = node498_r & ~pixel[709];
      node507_r = node506_l & pixel[187];
      node507_l = node506_l & ~pixel[187];
      node508 = node507_l;
      node509 = node507_r;
      node510 = node506_r;
      node511_r = node449_r & pixel[511];
      node511_l = node449_r & ~pixel[511];
      node512_r = node511_l & pixel[437];
      node512_l = node511_l & ~pixel[437];
      node513_r = node512_l & pixel[211];
      node513_l = node512_l & ~pixel[211];
      node514_r = node513_l & pixel[297];
      node514_l = node513_l & ~pixel[297];
      node515 = node514_l;
      node516_r = node514_r & pixel[349];
      node516_l = node514_r & ~pixel[349];
      node517 = node516_l;
      node518 = node516_r;
      node519_r = node513_r & pixel[409];
      node519_l = node513_r & ~pixel[409];
      node520_r = node519_l & pixel[203];
      node520_l = node519_l & ~pixel[203];
      node521 = node520_l;
      node522 = node520_r;
      node523 = node519_r;
      node524_r = node512_r & pixel[481];
      node524_l = node512_r & ~pixel[481];
      node525_r = node524_l & pixel[547];
      node525_l = node524_l & ~pixel[547];
      node526_r = node525_l & pixel[630];
      node526_l = node525_l & ~pixel[630];
      node527 = node526_l;
      node528 = node526_r;
      node529_r = node525_r & pixel[484];
      node529_l = node525_r & ~pixel[484];
      node530 = node529_l;
      node531 = node529_r;
      node532 = node524_r;
      node533_r = node511_r & pixel[408];
      node533_l = node511_r & ~pixel[408];
      node534_r = node533_l & pixel[431];
      node534_l = node533_l & ~pixel[431];
      node535_r = node534_l & pixel[743];
      node535_l = node534_l & ~pixel[743];
      node536_r = node535_l & pixel[145];
      node536_l = node535_l & ~pixel[145];
      node537 = node536_l;
      node538 = node536_r;
      node539 = node535_r;
      node540_r = node534_r & pixel[347];
      node540_l = node534_r & ~pixel[347];
      node541_r = node540_l & pixel[538];
      node541_l = node540_l & ~pixel[538];
      node542 = node541_l;
      node543 = node541_r;
      node544 = node540_r;
      node545_r = node533_r & pixel[443];
      node545_l = node533_r & ~pixel[443];
      node546_r = node545_l & pixel[234];
      node546_l = node545_l & ~pixel[234];
      node547_r = node546_l & pixel[302];
      node547_l = node546_l & ~pixel[302];
      node548 = node547_l;
      node549 = node547_r;
      node550_r = node546_r & pixel[346];
      node550_l = node546_r & ~pixel[346];
      node551 = node550_l;
      node552 = node550_r;
      node553_r = node545_r & pixel[285];
      node553_l = node545_r & ~pixel[285];
      node554_r = node553_l & pixel[179];
      node554_l = node553_l & ~pixel[179];
      node555 = node554_l;
      node556 = node554_r;
      node557_r = node553_r & pixel[264];
      node557_l = node553_r & ~pixel[264];
      node558 = node557_l;
      node559 = node557_r;
      node560_r = node448_r & pixel[514];
      node560_l = node448_r & ~pixel[514];
      node561_r = node560_l & pixel[353];
      node561_l = node560_l & ~pixel[353];
      node562_r = node561_l & pixel[241];
      node562_l = node561_l & ~pixel[241];
      node563_r = node562_l & pixel[438];
      node563_l = node562_l & ~pixel[438];
      node564_r = node563_l & pixel[151];
      node564_l = node563_l & ~pixel[151];
      node565_r = node564_l & pixel[186];
      node565_l = node564_l & ~pixel[186];
      node566 = node565_l;
      node567 = node565_r;
      node568_r = node564_r & pixel[434];
      node568_l = node564_r & ~pixel[434];
      node569 = node568_l;
      node570 = node568_r;
      node571_r = node563_r & pixel[490];
      node571_l = node563_r & ~pixel[490];
      node572_r = node571_l & pixel[468];
      node572_l = node571_l & ~pixel[468];
      node573 = node572_l;
      node574 = node572_r;
      node575_r = node571_r & pixel[400];
      node575_l = node571_r & ~pixel[400];
      node576 = node575_l;
      node577 = node575_r;
      node578_r = node562_r & pixel[413];
      node578_l = node562_r & ~pixel[413];
      node579_r = node578_l & pixel[216];
      node579_l = node578_l & ~pixel[216];
      node580_r = node579_l & pixel[567];
      node580_l = node579_l & ~pixel[567];
      node581 = node580_l;
      node582 = node580_r;
      node583_r = node579_r & pixel[265];
      node583_l = node579_r & ~pixel[265];
      node584 = node583_l;
      node585 = node583_r;
      node586_r = node578_r & pixel[568];
      node586_l = node578_r & ~pixel[568];
      node587_r = node586_l & pixel[329];
      node587_l = node586_l & ~pixel[329];
      node588 = node587_l;
      node589 = node587_r;
      node590_r = node586_r & pixel[602];
      node590_l = node586_r & ~pixel[602];
      node591 = node590_l;
      node592 = node590_r;
      node593_r = node561_r & pixel[606];
      node593_l = node561_r & ~pixel[606];
      node594_r = node593_l & pixel[460];
      node594_l = node593_l & ~pixel[460];
      node595_r = node594_l & pixel[550];
      node595_l = node594_l & ~pixel[550];
      node596_r = node595_l & pixel[152];
      node596_l = node595_l & ~pixel[152];
      node597 = node596_l;
      node598 = node596_r;
      node599_r = node595_r & pixel[717];
      node599_l = node595_r & ~pixel[717];
      node600 = node599_l;
      node601 = node599_r;
      node602_r = node594_r & pixel[238];
      node602_l = node594_r & ~pixel[238];
      node603_r = node602_l & pixel[68];
      node603_l = node602_l & ~pixel[68];
      node604 = node603_l;
      node605 = node603_r;
      node606_r = node602_r & pixel[232];
      node606_l = node602_r & ~pixel[232];
      node607 = node606_l;
      node608 = node606_r;
      node609_r = node593_r & pixel[374];
      node609_l = node593_r & ~pixel[374];
      node610_r = node609_l & pixel[719];
      node610_l = node609_l & ~pixel[719];
      node611_r = node610_l & pixel[466];
      node611_l = node610_l & ~pixel[466];
      node612 = node611_l;
      node613 = node611_r;
      node614_r = node610_r & pixel[486];
      node614_l = node610_r & ~pixel[486];
      node615 = node614_l;
      node616 = node614_r;
      node617_r = node609_r & pixel[189];
      node617_l = node609_r & ~pixel[189];
      node618_r = node617_l & pixel[497];
      node618_l = node617_l & ~pixel[497];
      node619 = node618_l;
      node620 = node618_r;
      node621_r = node617_r & pixel[488];
      node621_l = node617_r & ~pixel[488];
      node622 = node621_l;
      node623 = node621_r;
      node624_r = node560_r & pixel[657];
      node624_l = node560_r & ~pixel[657];
      node625_r = node624_l & pixel[653];
      node625_l = node624_l & ~pixel[653];
      node626_r = node625_l & pixel[528];
      node626_l = node625_l & ~pixel[528];
      node627_r = node626_l & pixel[243];
      node627_l = node626_l & ~pixel[243];
      node628_r = node627_l & pixel[382];
      node628_l = node627_l & ~pixel[382];
      node629 = node628_l;
      node630 = node628_r;
      node631_r = node627_r & pixel[387];
      node631_l = node627_r & ~pixel[387];
      node632 = node631_l;
      node633 = node631_r;
      node634_r = node626_r & pixel[453];
      node634_l = node626_r & ~pixel[453];
      node635_r = node634_l & pixel[232];
      node635_l = node634_l & ~pixel[232];
      node636 = node635_l;
      node637 = node635_r;
      node638_r = node634_r & pixel[285];
      node638_l = node634_r & ~pixel[285];
      node639 = node638_l;
      node640 = node638_r;
      node641_r = node625_r & pixel[513];
      node641_l = node625_r & ~pixel[513];
      node642_r = node641_l & pixel[459];
      node642_l = node641_l & ~pixel[459];
      node643_r = node642_l & pixel[218];
      node643_l = node642_l & ~pixel[218];
      node644 = node643_l;
      node645 = node643_r;
      node646_r = node642_r & pixel[190];
      node646_l = node642_r & ~pixel[190];
      node647 = node646_l;
      node648 = node646_r;
      node649_r = node641_r & pixel[705];
      node649_l = node641_r & ~pixel[705];
      node650_r = node649_l & pixel[433];
      node650_l = node649_l & ~pixel[433];
      node651 = node650_l;
      node652 = node650_r;
      node653_r = node649_r & pixel[319];
      node653_l = node649_r & ~pixel[319];
      node654 = node653_l;
      node655 = node653_r;
      node656_r = node624_r & pixel[569];
      node656_l = node624_r & ~pixel[569];
      node657_r = node656_l & pixel[324];
      node657_l = node656_l & ~pixel[324];
      node658_r = node657_l & pixel[370];
      node658_l = node657_l & ~pixel[370];
      node659_r = node658_l & pixel[354];
      node659_l = node658_l & ~pixel[354];
      node660 = node659_l;
      node661 = node659_r;
      node662 = node658_r;
      node663_r = node657_r & pixel[159];
      node663_l = node657_r & ~pixel[159];
      node664_r = node663_l & pixel[377];
      node664_l = node663_l & ~pixel[377];
      node665 = node664_l;
      node666 = node664_r;
      node667_r = node663_r & pixel[179];
      node667_l = node663_r & ~pixel[179];
      node668 = node667_l;
      node669 = node667_r;
      node670_r = node656_r & pixel[524];
      node670_l = node656_r & ~pixel[524];
      node671_r = node670_l & pixel[461];
      node671_l = node670_l & ~pixel[461];
      node672_r = node671_l & pixel[219];
      node672_l = node671_l & ~pixel[219];
      node673 = node672_l;
      node674 = node672_r;
      node675_r = node671_r & pixel[609];
      node675_l = node671_r & ~pixel[609];
      node676 = node675_l;
      node677 = node675_r;
      node678_r = node670_r & pixel[232];
      node678_l = node670_r & ~pixel[232];
      node679_r = node678_l & pixel[191];
      node679_l = node678_l & ~pixel[191];
      node680 = node679_l;
      node681 = node679_r;
      node682_r = node678_r & pixel[488];
      node682_l = node678_r & ~pixel[488];
      node683 = node682_l;
      node684 = node682_r;
      node685_r = node447_r & pixel[497];
      node685_l = node447_r & ~pixel[497];
      node686_r = node685_l & pixel[213];
      node686_l = node685_l & ~pixel[213];
      node687_r = node686_l & pixel[245];
      node687_l = node686_l & ~pixel[245];
      node688_r = node687_l & pixel[125];
      node688_l = node687_l & ~pixel[125];
      node689_r = node688_l & pixel[261];
      node689_l = node688_l & ~pixel[261];
      node690_r = node689_l & pixel[244];
      node690_l = node689_l & ~pixel[244];
      node691_r = node690_l & pixel[238];
      node691_l = node690_l & ~pixel[238];
      node692 = node691_l;
      node693 = node691_r;
      node694_r = node690_r & pixel[71];
      node694_l = node690_r & ~pixel[71];
      node695 = node694_l;
      node696 = node694_r;
      node697_r = node689_r & pixel[297];
      node697_l = node689_r & ~pixel[297];
      node698_r = node697_l & pixel[490];
      node698_l = node697_l & ~pixel[490];
      node699 = node698_l;
      node700 = node698_r;
      node701_r = node697_r & pixel[236];
      node701_l = node697_r & ~pixel[236];
      node702 = node701_l;
      node703 = node701_r;
      node704_r = node688_r & pixel[633];
      node704_l = node688_r & ~pixel[633];
      node705_r = node704_l & pixel[302];
      node705_l = node704_l & ~pixel[302];
      node706_r = node705_l & pixel[187];
      node706_l = node705_l & ~pixel[187];
      node707 = node706_l;
      node708 = node706_r;
      node709_r = node705_r & pixel[522];
      node709_l = node705_r & ~pixel[522];
      node710 = node709_l;
      node711 = node709_r;
      node712_r = node704_r & pixel[345];
      node712_l = node704_r & ~pixel[345];
      node713_r = node712_l & pixel[544];
      node713_l = node712_l & ~pixel[544];
      node714 = node713_l;
      node715 = node713_r;
      node716_r = node712_r & pixel[427];
      node716_l = node712_r & ~pixel[427];
      node717 = node716_l;
      node718 = node716_r;
      node719_r = node687_r & pixel[277];
      node719_l = node687_r & ~pixel[277];
      node720_r = node719_l & pixel[327];
      node720_l = node719_l & ~pixel[327];
      node721_r = node720_l & pixel[454];
      node721_l = node720_l & ~pixel[454];
      node722_r = node721_l & pixel[543];
      node722_l = node721_l & ~pixel[543];
      node723 = node722_l;
      node724 = node722_r;
      node725_r = node721_r & pixel[438];
      node725_l = node721_r & ~pixel[438];
      node726 = node725_l;
      node727 = node725_r;
      node728_r = node720_r & pixel[239];
      node728_l = node720_r & ~pixel[239];
      node729_r = node728_l & pixel[268];
      node729_l = node728_l & ~pixel[268];
      node730 = node729_l;
      node731 = node729_r;
      node732_r = node728_r & pixel[431];
      node732_l = node728_r & ~pixel[431];
      node733 = node732_l;
      node734 = node732_r;
      node735_r = node719_r & pixel[352];
      node735_l = node719_r & ~pixel[352];
      node736_r = node735_l & pixel[411];
      node736_l = node735_l & ~pixel[411];
      node737 = node736_l;
      node738 = node736_r;
      node739_r = node735_r & pixel[384];
      node739_l = node735_r & ~pixel[384];
      node740_r = node739_l & pixel[379];
      node740_l = node739_l & ~pixel[379];
      node741 = node740_l;
      node742 = node740_r;
      node743_r = node739_r & pixel[232];
      node743_l = node739_r & ~pixel[232];
      node744 = node743_l;
      node745 = node743_r;
      node746_r = node686_r & pixel[408];
      node746_l = node686_r & ~pixel[408];
      node747_r = node746_l & pixel[467];
      node747_l = node746_l & ~pixel[467];
      node748_r = node747_l & pixel[438];
      node748_l = node747_l & ~pixel[438];
      node749_r = node748_l & pixel[353];
      node749_l = node748_l & ~pixel[353];
      node750_r = node749_l & pixel[527];
      node750_l = node749_l & ~pixel[527];
      node751 = node750_l;
      node752 = node750_r;
      node753_r = node749_r & pixel[461];
      node753_l = node749_r & ~pixel[461];
      node754 = node753_l;
      node755 = node753_r;
      node756_r = node748_r & pixel[490];
      node756_l = node748_r & ~pixel[490];
      node757_r = node756_l & pixel[349];
      node757_l = node756_l & ~pixel[349];
      node758 = node757_l;
      node759 = node757_r;
      node760_r = node756_r & pixel[354];
      node760_l = node756_r & ~pixel[354];
      node761 = node760_l;
      node762 = node760_r;
      node763_r = node747_r & pixel[347];
      node763_l = node747_r & ~pixel[347];
      node764_r = node763_l & pixel[555];
      node764_l = node763_l & ~pixel[555];
      node765_r = node764_l & pixel[239];
      node765_l = node764_l & ~pixel[239];
      node766 = node765_l;
      node767 = node765_r;
      node768 = node764_r;
      node769_r = node763_r & pixel[412];
      node769_l = node763_r & ~pixel[412];
      node770_r = node769_l & pixel[99];
      node770_l = node769_l & ~pixel[99];
      node771 = node770_l;
      node772 = node770_r;
      node773_r = node769_r & pixel[321];
      node773_l = node769_r & ~pixel[321];
      node774 = node773_l;
      node775 = node773_r;
      node776_r = node746_r & pixel[325];
      node776_l = node746_r & ~pixel[325];
      node777_r = node776_l & pixel[192];
      node777_l = node776_l & ~pixel[192];
      node778_r = node777_l & pixel[326];
      node778_l = node777_l & ~pixel[326];
      node779_r = node778_l & pixel[517];
      node779_l = node778_l & ~pixel[517];
      node780 = node779_l;
      node781 = node779_r;
      node782_r = node778_r & pixel[611];
      node782_l = node778_r & ~pixel[611];
      node783 = node782_l;
      node784 = node782_r;
      node785_r = node777_r & pixel[358];
      node785_l = node777_r & ~pixel[358];
      node786_r = node785_l & pixel[576];
      node786_l = node785_l & ~pixel[576];
      node787 = node786_l;
      node788 = node786_r;
      node789_r = node785_r & pixel[462];
      node789_l = node785_r & ~pixel[462];
      node790 = node789_l;
      node791 = node789_r;
      node792_r = node776_r & pixel[622];
      node792_l = node776_r & ~pixel[622];
      node793_r = node792_l & pixel[710];
      node793_l = node792_l & ~pixel[710];
      node794_r = node793_l & pixel[598];
      node794_l = node793_l & ~pixel[598];
      node795 = node794_l;
      node796 = node794_r;
      node797_r = node793_r & pixel[233];
      node797_l = node793_r & ~pixel[233];
      node798 = node797_l;
      node799 = node797_r;
      node800_r = node792_r & pixel[517];
      node800_l = node792_r & ~pixel[517];
      node801_r = node800_l & pixel[607];
      node801_l = node800_l & ~pixel[607];
      node802 = node801_l;
      node803 = node801_r;
      node804_r = node800_r & pixel[212];
      node804_l = node800_r & ~pixel[212];
      node805 = node804_l;
      node806 = node804_r;
      node807_r = node685_r & pixel[241];
      node807_l = node685_r & ~pixel[241];
      node808_r = node807_l & pixel[95];
      node808_l = node807_l & ~pixel[95];
      node809_r = node808_l & pixel[543];
      node809_l = node808_l & ~pixel[543];
      node810_r = node809_l & pixel[492];
      node810_l = node809_l & ~pixel[492];
      node811_r = node810_l & pixel[213];
      node811_l = node810_l & ~pixel[213];
      node812_r = node811_l & pixel[686];
      node812_l = node811_l & ~pixel[686];
      node813 = node812_l;
      node814 = node812_r;
      node815_r = node811_r & pixel[522];
      node815_l = node811_r & ~pixel[522];
      node816 = node815_l;
      node817 = node815_r;
      node818_r = node810_r & pixel[218];
      node818_l = node810_r & ~pixel[218];
      node819_r = node818_l & pixel[321];
      node819_l = node818_l & ~pixel[321];
      node820 = node819_l;
      node821 = node819_r;
      node822_r = node818_r & pixel[624];
      node822_l = node818_r & ~pixel[624];
      node823 = node822_l;
      node824 = node822_r;
      node825_r = node809_r & pixel[99];
      node825_l = node809_r & ~pixel[99];
      node826_r = node825_l & pixel[124];
      node826_l = node825_l & ~pixel[124];
      node827_r = node826_l & pixel[327];
      node827_l = node826_l & ~pixel[327];
      node828 = node827_l;
      node829 = node827_r;
      node830_r = node826_r & pixel[566];
      node830_l = node826_r & ~pixel[566];
      node831 = node830_l;
      node832 = node830_r;
      node833 = node825_r;
      node834_r = node808_r & pixel[543];
      node834_l = node808_r & ~pixel[543];
      node835_r = node834_l & pixel[126];
      node835_l = node834_l & ~pixel[126];
      node836 = node835_l;
      node837 = node835_r;
      node838_r = node834_r & pixel[234];
      node838_l = node834_r & ~pixel[234];
      node839_r = node838_l & pixel[96];
      node839_l = node838_l & ~pixel[96];
      node840 = node839_l;
      node841 = node839_r;
      node842_r = node838_r & pixel[264];
      node842_l = node838_r & ~pixel[264];
      node843 = node842_l;
      node844_r = node842_r & pixel[631];
      node844_l = node842_r & ~pixel[631];
      node845 = node844_l;
      node846 = node844_r;
      node847_r = node807_r & pixel[598];
      node847_l = node807_r & ~pixel[598];
      node848_r = node847_l & pixel[552];
      node848_l = node847_l & ~pixel[552];
      node849_r = node848_l & pixel[187];
      node849_l = node848_l & ~pixel[187];
      node850_r = node849_l & pixel[266];
      node850_l = node849_l & ~pixel[266];
      node851_r = node850_l & pixel[467];
      node851_l = node850_l & ~pixel[467];
      node852 = node851_l;
      node853 = node851_r;
      node854_r = node850_r & pixel[541];
      node854_l = node850_r & ~pixel[541];
      node855 = node854_l;
      node856 = node854_r;
      node857_r = node849_r & pixel[464];
      node857_l = node849_r & ~pixel[464];
      node858_r = node857_l & pixel[541];
      node858_l = node857_l & ~pixel[541];
      node859 = node858_l;
      node860 = node858_r;
      node861_r = node857_r & pixel[547];
      node861_l = node857_r & ~pixel[547];
      node862 = node861_l;
      node863 = node861_r;
      node864_r = node848_r & pixel[655];
      node864_l = node848_r & ~pixel[655];
      node865_r = node864_l & pixel[239];
      node865_l = node864_l & ~pixel[239];
      node866_r = node865_l & pixel[456];
      node866_l = node865_l & ~pixel[456];
      node867 = node866_l;
      node868 = node866_r;
      node869_r = node865_r & pixel[666];
      node869_l = node865_r & ~pixel[666];
      node870 = node869_l;
      node871 = node869_r;
      node872_r = node864_r & pixel[326];
      node872_l = node864_r & ~pixel[326];
      node873_r = node872_l & pixel[538];
      node873_l = node872_l & ~pixel[538];
      node874 = node873_l;
      node875 = node873_r;
      node876_r = node872_r & pixel[178];
      node876_l = node872_r & ~pixel[178];
      node877 = node876_l;
      node878 = node876_r;
      node879_r = node847_r & pixel[379];
      node879_l = node847_r & ~pixel[379];
      node880_r = node879_l & pixel[289];
      node880_l = node879_l & ~pixel[289];
      node881_r = node880_l & pixel[217];
      node881_l = node880_l & ~pixel[217];
      node882_r = node881_l & pixel[381];
      node882_l = node881_l & ~pixel[381];
      node883 = node882_l;
      node884 = node882_r;
      node885_r = node881_r & pixel[318];
      node885_l = node881_r & ~pixel[318];
      node886 = node885_l;
      node887 = node885_r;
      node888_r = node880_r & pixel[405];
      node888_l = node880_r & ~pixel[405];
      node889_r = node888_l & pixel[249];
      node889_l = node888_l & ~pixel[249];
      node890 = node889_l;
      node891 = node889_r;
      node892_r = node888_r & pixel[302];
      node892_l = node888_r & ~pixel[302];
      node893 = node892_l;
      node894 = node892_r;
      node895_r = node879_r & pixel[630];
      node895_l = node879_r & ~pixel[630];
      node896_r = node895_l & pixel[373];
      node896_l = node895_l & ~pixel[373];
      node897_r = node896_l & pixel[509];
      node897_l = node896_l & ~pixel[509];
      node898 = node897_l;
      node899 = node897_r;
      node900_r = node896_r & pixel[239];
      node900_l = node896_r & ~pixel[239];
      node901 = node900_l;
      node902 = node900_r;
      node903_r = node895_r & pixel[455];
      node903_l = node895_r & ~pixel[455];
      node904_r = node903_l & pixel[355];
      node904_l = node903_l & ~pixel[355];
      node905 = node904_l;
      node906 = node904_r;
      node907_r = node903_r & pixel[486];
      node907_l = node903_r & ~pixel[486];
      node908 = node907_l;
      node909 = node907_r;
      node910_r = node0_r & pixel[488];
      node910_l = node0_r & ~pixel[488];
      node911_r = node910_l & pixel[317];
      node911_l = node910_l & ~pixel[317];
      node912_r = node911_l & pixel[270];
      node912_l = node911_l & ~pixel[270];
      node913_r = node912_l & pixel[655];
      node913_l = node912_l & ~pixel[655];
      node914_r = node913_l & pixel[430];
      node914_l = node913_l & ~pixel[430];
      node915_r = node914_l & pixel[493];
      node915_l = node914_l & ~pixel[493];
      node916_r = node915_l & pixel[625];
      node916_l = node915_l & ~pixel[625];
      node917_r = node916_l & pixel[205];
      node917_l = node916_l & ~pixel[205];
      node918_r = node917_l & pixel[599];
      node918_l = node917_l & ~pixel[599];
      node919 = node918_l;
      node920 = node918_r;
      node921_r = node917_r & pixel[375];
      node921_l = node917_r & ~pixel[375];
      node922 = node921_l;
      node923 = node921_r;
      node924_r = node916_r & pixel[126];
      node924_l = node916_r & ~pixel[126];
      node925_r = node924_l & pixel[398];
      node925_l = node924_l & ~pixel[398];
      node926 = node925_l;
      node927 = node925_r;
      node928_r = node924_r & pixel[187];
      node928_l = node924_r & ~pixel[187];
      node929 = node928_l;
      node930 = node928_r;
      node931_r = node915_r & pixel[327];
      node931_l = node915_r & ~pixel[327];
      node932_r = node931_l & pixel[295];
      node932_l = node931_l & ~pixel[295];
      node933_r = node932_l & pixel[341];
      node933_l = node932_l & ~pixel[341];
      node934 = node933_l;
      node935 = node933_r;
      node936_r = node932_r & pixel[518];
      node936_l = node932_r & ~pixel[518];
      node937 = node936_l;
      node938 = node936_r;
      node939_r = node931_r & pixel[426];
      node939_l = node931_r & ~pixel[426];
      node940_r = node939_l & pixel[408];
      node940_l = node939_l & ~pixel[408];
      node941 = node940_l;
      node942 = node940_r;
      node943 = node939_r;
      node944_r = node914_r & pixel[245];
      node944_l = node914_r & ~pixel[245];
      node945_r = node944_l & pixel[528];
      node945_l = node944_l & ~pixel[528];
      node946_r = node945_l & pixel[129];
      node946_l = node945_l & ~pixel[129];
      node947_r = node946_l & pixel[179];
      node947_l = node946_l & ~pixel[179];
      node948 = node947_l;
      node949 = node947_r;
      node950_r = node946_r & pixel[179];
      node950_l = node946_r & ~pixel[179];
      node951 = node950_l;
      node952 = node950_r;
      node953_r = node945_r & pixel[512];
      node953_l = node945_r & ~pixel[512];
      node954_r = node953_l & pixel[243];
      node954_l = node953_l & ~pixel[243];
      node955 = node954_l;
      node956 = node954_r;
      node957_r = node953_r & pixel[263];
      node957_l = node953_r & ~pixel[263];
      node958 = node957_l;
      node959 = node957_r;
      node960_r = node944_r & pixel[349];
      node960_l = node944_r & ~pixel[349];
      node961_r = node960_l & pixel[346];
      node961_l = node960_l & ~pixel[346];
      node962_r = node961_l & pixel[481];
      node962_l = node961_l & ~pixel[481];
      node963 = node962_l;
      node964 = node962_r;
      node965 = node961_r;
      node966_r = node960_r & pixel[324];
      node966_l = node960_r & ~pixel[324];
      node967_r = node966_l & pixel[293];
      node967_l = node966_l & ~pixel[293];
      node968 = node967_l;
      node969 = node967_r;
      node970 = node966_r;
      node971_r = node913_r & pixel[216];
      node971_l = node913_r & ~pixel[216];
      node972_r = node971_l & pixel[264];
      node972_l = node971_l & ~pixel[264];
      node973_r = node972_l & pixel[376];
      node973_l = node972_l & ~pixel[376];
      node974_r = node973_l & pixel[522];
      node974_l = node973_l & ~pixel[522];
      node975_r = node974_l & pixel[573];
      node975_l = node974_l & ~pixel[573];
      node976 = node975_l;
      node977 = node975_r;
      node978_r = node974_r & pixel[517];
      node978_l = node974_r & ~pixel[517];
      node979 = node978_l;
      node980 = node978_r;
      node981_r = node973_r & pixel[268];
      node981_l = node973_r & ~pixel[268];
      node982_r = node981_l & pixel[290];
      node982_l = node981_l & ~pixel[290];
      node983 = node982_l;
      node984 = node982_r;
      node985_r = node981_r & pixel[163];
      node985_l = node981_r & ~pixel[163];
      node986 = node985_l;
      node987 = node985_r;
      node988_r = node972_r & pixel[159];
      node988_l = node972_r & ~pixel[159];
      node989_r = node988_l & pixel[212];
      node989_l = node988_l & ~pixel[212];
      node990_r = node989_l & pixel[490];
      node990_l = node989_l & ~pixel[490];
      node991 = node990_l;
      node992 = node990_r;
      node993_r = node989_r & pixel[467];
      node993_l = node989_r & ~pixel[467];
      node994 = node993_l;
      node995 = node993_r;
      node996_r = node988_r & pixel[273];
      node996_l = node988_r & ~pixel[273];
      node997_r = node996_l & pixel[268];
      node997_l = node996_l & ~pixel[268];
      node998 = node997_l;
      node999 = node997_r;
      node1000_r = node996_r & pixel[375];
      node1000_l = node996_r & ~pixel[375];
      node1001 = node1000_l;
      node1002 = node1000_r;
      node1003_r = node971_r & pixel[414];
      node1003_l = node971_r & ~pixel[414];
      node1004_r = node1003_l & pixel[379];
      node1004_l = node1003_l & ~pixel[379];
      node1005_r = node1004_l & pixel[688];
      node1005_l = node1004_l & ~pixel[688];
      node1006_r = node1005_l & pixel[536];
      node1006_l = node1005_l & ~pixel[536];
      node1007 = node1006_l;
      node1008 = node1006_r;
      node1009_r = node1005_r & pixel[236];
      node1009_l = node1005_r & ~pixel[236];
      node1010 = node1009_l;
      node1011 = node1009_r;
      node1012_r = node1004_r & pixel[328];
      node1012_l = node1004_r & ~pixel[328];
      node1013_r = node1012_l & pixel[273];
      node1013_l = node1012_l & ~pixel[273];
      node1014 = node1013_l;
      node1015 = node1013_r;
      node1016_r = node1012_r & pixel[549];
      node1016_l = node1012_r & ~pixel[549];
      node1017 = node1016_l;
      node1018 = node1016_r;
      node1019_r = node1003_r & pixel[563];
      node1019_l = node1003_r & ~pixel[563];
      node1020_r = node1019_l & pixel[324];
      node1020_l = node1019_l & ~pixel[324];
      node1021_r = node1020_l & pixel[354];
      node1021_l = node1020_l & ~pixel[354];
      node1022 = node1021_l;
      node1023 = node1021_r;
      node1024_r = node1020_r & pixel[121];
      node1024_l = node1020_r & ~pixel[121];
      node1025 = node1024_l;
      node1026 = node1024_r;
      node1027 = node1019_r;
      node1028_r = node912_r & pixel[323];
      node1028_l = node912_r & ~pixel[323];
      node1029_r = node1028_l & pixel[492];
      node1029_l = node1028_l & ~pixel[492];
      node1030_r = node1029_l & pixel[408];
      node1030_l = node1029_l & ~pixel[408];
      node1031_r = node1030_l & pixel[96];
      node1031_l = node1030_l & ~pixel[96];
      node1032_r = node1031_l & pixel[463];
      node1032_l = node1031_l & ~pixel[463];
      node1033_r = node1032_l & pixel[518];
      node1033_l = node1032_l & ~pixel[518];
      node1034 = node1033_l;
      node1035 = node1033_r;
      node1036_r = node1032_r & pixel[120];
      node1036_l = node1032_r & ~pixel[120];
      node1037 = node1036_l;
      node1038 = node1036_r;
      node1039_r = node1031_r & pixel[385];
      node1039_l = node1031_r & ~pixel[385];
      node1040 = node1039_l;
      node1041 = node1039_r;
      node1042_r = node1030_r & pixel[632];
      node1042_l = node1030_r & ~pixel[632];
      node1043_r = node1042_l & pixel[571];
      node1043_l = node1042_l & ~pixel[571];
      node1044_r = node1043_l & pixel[372];
      node1044_l = node1043_l & ~pixel[372];
      node1045 = node1044_l;
      node1046 = node1044_r;
      node1047_r = node1043_r & pixel[123];
      node1047_l = node1043_r & ~pixel[123];
      node1048 = node1047_l;
      node1049 = node1047_r;
      node1050_r = node1042_r & pixel[427];
      node1050_l = node1042_r & ~pixel[427];
      node1051_r = node1050_l & pixel[244];
      node1051_l = node1050_l & ~pixel[244];
      node1052 = node1051_l;
      node1053 = node1051_r;
      node1054_r = node1050_r & pixel[341];
      node1054_l = node1050_r & ~pixel[341];
      node1055 = node1054_l;
      node1056 = node1054_r;
      node1057_r = node1029_r & pixel[462];
      node1057_l = node1029_r & ~pixel[462];
      node1058_r = node1057_l & pixel[176];
      node1058_l = node1057_l & ~pixel[176];
      node1059_r = node1058_l & pixel[293];
      node1059_l = node1058_l & ~pixel[293];
      node1060_r = node1059_l & pixel[569];
      node1060_l = node1059_l & ~pixel[569];
      node1061 = node1060_l;
      node1062 = node1060_r;
      node1063_r = node1059_r & pixel[513];
      node1063_l = node1059_r & ~pixel[513];
      node1064 = node1063_l;
      node1065 = node1063_r;
      node1066_r = node1058_r & pixel[185];
      node1066_l = node1058_r & ~pixel[185];
      node1067_r = node1066_l & pixel[605];
      node1067_l = node1066_l & ~pixel[605];
      node1068 = node1067_l;
      node1069 = node1067_r;
      node1070_r = node1066_r & pixel[572];
      node1070_l = node1066_r & ~pixel[572];
      node1071 = node1070_l;
      node1072 = node1070_r;
      node1073_r = node1057_r & pixel[455];
      node1073_l = node1057_r & ~pixel[455];
      node1074_r = node1073_l & pixel[512];
      node1074_l = node1073_l & ~pixel[512];
      node1075_r = node1074_l & pixel[571];
      node1075_l = node1074_l & ~pixel[571];
      node1076 = node1075_l;
      node1077 = node1075_r;
      node1078_r = node1074_r & pixel[379];
      node1078_l = node1074_r & ~pixel[379];
      node1079 = node1078_l;
      node1080 = node1078_r;
      node1081_r = node1073_r & pixel[429];
      node1081_l = node1073_r & ~pixel[429];
      node1082_r = node1081_l & pixel[301];
      node1082_l = node1081_l & ~pixel[301];
      node1083 = node1082_l;
      node1084 = node1082_r;
      node1085_r = node1081_r & pixel[293];
      node1085_l = node1081_r & ~pixel[293];
      node1086 = node1085_l;
      node1087 = node1085_r;
      node1088_r = node1028_r & pixel[654];
      node1088_l = node1028_r & ~pixel[654];
      node1089_r = node1088_l & pixel[485];
      node1089_l = node1088_l & ~pixel[485];
      node1090_r = node1089_l & pixel[350];
      node1090_l = node1089_l & ~pixel[350];
      node1091_r = node1090_l & pixel[353];
      node1091_l = node1090_l & ~pixel[353];
      node1092_r = node1091_l & pixel[160];
      node1092_l = node1091_l & ~pixel[160];
      node1093 = node1092_l;
      node1094 = node1092_r;
      node1095_r = node1091_r & pixel[97];
      node1095_l = node1091_r & ~pixel[97];
      node1096 = node1095_l;
      node1097 = node1095_r;
      node1098_r = node1090_r & pixel[487];
      node1098_l = node1090_r & ~pixel[487];
      node1099_r = node1098_l & pixel[666];
      node1099_l = node1098_l & ~pixel[666];
      node1100 = node1099_l;
      node1101 = node1099_r;
      node1102_r = node1098_r & pixel[517];
      node1102_l = node1098_r & ~pixel[517];
      node1103 = node1102_l;
      node1104 = node1102_r;
      node1105_r = node1089_r & pixel[431];
      node1105_l = node1089_r & ~pixel[431];
      node1106_r = node1105_l & pixel[318];
      node1106_l = node1105_l & ~pixel[318];
      node1107_r = node1106_l & pixel[509];
      node1107_l = node1106_l & ~pixel[509];
      node1108 = node1107_l;
      node1109 = node1107_r;
      node1110_r = node1106_r & pixel[661];
      node1110_l = node1106_r & ~pixel[661];
      node1111 = node1110_l;
      node1112 = node1110_r;
      node1113_r = node1105_r & pixel[656];
      node1113_l = node1105_r & ~pixel[656];
      node1114_r = node1113_l & pixel[631];
      node1114_l = node1113_l & ~pixel[631];
      node1115 = node1114_l;
      node1116 = node1114_r;
      node1117_r = node1113_r & pixel[177];
      node1117_l = node1113_r & ~pixel[177];
      node1118 = node1117_l;
      node1119 = node1117_r;
      node1120_r = node1088_r & pixel[458];
      node1120_l = node1088_r & ~pixel[458];
      node1121_r = node1120_l & pixel[292];
      node1121_l = node1120_l & ~pixel[292];
      node1122_r = node1121_l & pixel[331];
      node1122_l = node1121_l & ~pixel[331];
      node1123_r = node1122_l & pixel[156];
      node1123_l = node1122_l & ~pixel[156];
      node1124 = node1123_l;
      node1125 = node1123_r;
      node1126_r = node1122_r & pixel[188];
      node1126_l = node1122_r & ~pixel[188];
      node1127 = node1126_l;
      node1128 = node1126_r;
      node1129_r = node1121_r & pixel[438];
      node1129_l = node1121_r & ~pixel[438];
      node1130_r = node1129_l & pixel[176];
      node1130_l = node1129_l & ~pixel[176];
      node1131 = node1130_l;
      node1132 = node1130_r;
      node1133_r = node1129_r & pixel[350];
      node1133_l = node1129_r & ~pixel[350];
      node1134 = node1133_l;
      node1135 = node1133_r;
      node1136_r = node1120_r & pixel[206];
      node1136_l = node1120_r & ~pixel[206];
      node1137_r = node1136_l & pixel[384];
      node1137_l = node1136_l & ~pixel[384];
      node1138_r = node1137_l & pixel[484];
      node1138_l = node1137_l & ~pixel[484];
      node1139 = node1138_l;
      node1140 = node1138_r;
      node1141_r = node1137_r & pixel[433];
      node1141_l = node1137_r & ~pixel[433];
      node1142 = node1141_l;
      node1143 = node1141_r;
      node1144_r = node1136_r & pixel[541];
      node1144_l = node1136_r & ~pixel[541];
      node1145_r = node1144_l & pixel[540];
      node1145_l = node1144_l & ~pixel[540];
      node1146 = node1145_l;
      node1147 = node1145_r;
      node1148_r = node1144_r & pixel[523];
      node1148_l = node1144_r & ~pixel[523];
      node1149 = node1148_l;
      node1150 = node1148_r;
      node1151_r = node911_r & pixel[409];
      node1151_l = node911_r & ~pixel[409];
      node1152_r = node1151_l & pixel[413];
      node1152_l = node1151_l & ~pixel[413];
      node1153_r = node1152_l & pixel[387];
      node1153_l = node1152_l & ~pixel[387];
      node1154_r = node1153_l & pixel[456];
      node1154_l = node1153_l & ~pixel[456];
      node1155_r = node1154_l & pixel[187];
      node1155_l = node1154_l & ~pixel[187];
      node1156_r = node1155_l & pixel[515];
      node1156_l = node1155_l & ~pixel[515];
      node1157_r = node1156_l & pixel[240];
      node1157_l = node1156_l & ~pixel[240];
      node1158 = node1157_l;
      node1159 = node1157_r;
      node1160_r = node1156_r & pixel[519];
      node1160_l = node1156_r & ~pixel[519];
      node1161 = node1160_l;
      node1162 = node1160_r;
      node1163_r = node1155_r & pixel[326];
      node1163_l = node1155_r & ~pixel[326];
      node1164_r = node1163_l & pixel[294];
      node1164_l = node1163_l & ~pixel[294];
      node1165 = node1164_l;
      node1166 = node1164_r;
      node1167_r = node1163_r & pixel[486];
      node1167_l = node1163_r & ~pixel[486];
      node1168 = node1167_l;
      node1169 = node1167_r;
      node1170_r = node1154_r & pixel[435];
      node1170_l = node1154_r & ~pixel[435];
      node1171_r = node1170_l & pixel[490];
      node1171_l = node1170_l & ~pixel[490];
      node1172_r = node1171_l & pixel[271];
      node1172_l = node1171_l & ~pixel[271];
      node1173 = node1172_l;
      node1174 = node1172_r;
      node1175_r = node1171_r & pixel[373];
      node1175_l = node1171_r & ~pixel[373];
      node1176 = node1175_l;
      node1177 = node1175_r;
      node1178_r = node1170_r & pixel[438];
      node1178_l = node1170_r & ~pixel[438];
      node1179_r = node1178_l & pixel[296];
      node1179_l = node1178_l & ~pixel[296];
      node1180 = node1179_l;
      node1181 = node1179_r;
      node1182_r = node1178_r & pixel[100];
      node1182_l = node1178_r & ~pixel[100];
      node1183 = node1182_l;
      node1184 = node1182_r;
      node1185_r = node1153_r & pixel[147];
      node1185_l = node1153_r & ~pixel[147];
      node1186_r = node1185_l & pixel[382];
      node1186_l = node1185_l & ~pixel[382];
      node1187_r = node1186_l & pixel[302];
      node1187_l = node1186_l & ~pixel[302];
      node1188_r = node1187_l & pixel[472];
      node1188_l = node1187_l & ~pixel[472];
      node1189 = node1188_l;
      node1190 = node1188_r;
      node1191 = node1187_r;
      node1192_r = node1186_r & pixel[275];
      node1192_l = node1186_r & ~pixel[275];
      node1193_r = node1192_l & pixel[231];
      node1193_l = node1192_l & ~pixel[231];
      node1194 = node1193_l;
      node1195 = node1193_r;
      node1196 = node1192_r;
      node1197_r = node1185_r & pixel[331];
      node1197_l = node1185_r & ~pixel[331];
      node1198 = node1197_l;
      node1199_r = node1197_r & pixel[295];
      node1199_l = node1197_r & ~pixel[295];
      node1200 = node1199_l;
      node1201 = node1199_r;
      node1202_r = node1152_r & pixel[382];
      node1202_l = node1152_r & ~pixel[382];
      node1203_r = node1202_l & pixel[406];
      node1203_l = node1202_l & ~pixel[406];
      node1204_r = node1203_l & pixel[400];
      node1204_l = node1203_l & ~pixel[400];
      node1205_r = node1204_l & pixel[353];
      node1205_l = node1204_l & ~pixel[353];
      node1206_r = node1205_l & pixel[119];
      node1206_l = node1205_l & ~pixel[119];
      node1207 = node1206_l;
      node1208 = node1206_r;
      node1209_r = node1205_r & pixel[600];
      node1209_l = node1205_r & ~pixel[600];
      node1210 = node1209_l;
      node1211 = node1209_r;
      node1212_r = node1204_r & pixel[329];
      node1212_l = node1204_r & ~pixel[329];
      node1213_r = node1212_l & pixel[605];
      node1213_l = node1212_l & ~pixel[605];
      node1214 = node1213_l;
      node1215 = node1213_r;
      node1216_r = node1212_r & pixel[378];
      node1216_l = node1212_r & ~pixel[378];
      node1217 = node1216_l;
      node1218 = node1216_r;
      node1219_r = node1203_r & pixel[263];
      node1219_l = node1203_r & ~pixel[263];
      node1220_r = node1219_l & pixel[491];
      node1220_l = node1219_l & ~pixel[491];
      node1221 = node1220_l;
      node1222 = node1220_r;
      node1223_r = node1219_r & pixel[605];
      node1223_l = node1219_r & ~pixel[605];
      node1224_r = node1223_l & pixel[466];
      node1224_l = node1223_l & ~pixel[466];
      node1225 = node1224_l;
      node1226 = node1224_r;
      node1227_r = node1223_r & pixel[358];
      node1227_l = node1223_r & ~pixel[358];
      node1228 = node1227_l;
      node1229 = node1227_r;
      node1230_r = node1202_r & pixel[325];
      node1230_l = node1202_r & ~pixel[325];
      node1231_r = node1230_l & pixel[380];
      node1231_l = node1230_l & ~pixel[380];
      node1232_r = node1231_l & pixel[596];
      node1232_l = node1231_l & ~pixel[596];
      node1233_r = node1232_l & pixel[691];
      node1233_l = node1232_l & ~pixel[691];
      node1234 = node1233_l;
      node1235 = node1233_r;
      node1236 = node1232_r;
      node1237_r = node1231_r & pixel[633];
      node1237_l = node1231_r & ~pixel[633];
      node1238 = node1237_l;
      node1239_r = node1237_r & pixel[397];
      node1239_l = node1237_r & ~pixel[397];
      node1240 = node1239_l;
      node1241 = node1239_r;
      node1242_r = node1230_r & pixel[427];
      node1242_l = node1230_r & ~pixel[427];
      node1243_r = node1242_l & pixel[287];
      node1243_l = node1242_l & ~pixel[287];
      node1244_r = node1243_l & pixel[263];
      node1244_l = node1243_l & ~pixel[263];
      node1245 = node1244_l;
      node1246 = node1244_r;
      node1247_r = node1243_r & pixel[469];
      node1247_l = node1243_r & ~pixel[469];
      node1248 = node1247_l;
      node1249 = node1247_r;
      node1250_r = node1242_r & pixel[377];
      node1250_l = node1242_r & ~pixel[377];
      node1251_r = node1250_l & pixel[262];
      node1251_l = node1250_l & ~pixel[262];
      node1252 = node1251_l;
      node1253 = node1251_r;
      node1254_r = node1250_r & pixel[484];
      node1254_l = node1250_r & ~pixel[484];
      node1255 = node1254_l;
      node1256 = node1254_r;
      node1257_r = node1151_r & pixel[455];
      node1257_l = node1151_r & ~pixel[455];
      node1258_r = node1257_l & pixel[289];
      node1258_l = node1257_l & ~pixel[289];
      node1259_r = node1258_l & pixel[513];
      node1259_l = node1258_l & ~pixel[513];
      node1260_r = node1259_l & pixel[151];
      node1260_l = node1259_l & ~pixel[151];
      node1261_r = node1260_l & pixel[507];
      node1261_l = node1260_l & ~pixel[507];
      node1262_r = node1261_l & pixel[466];
      node1262_l = node1261_l & ~pixel[466];
      node1263 = node1262_l;
      node1264 = node1262_r;
      node1265 = node1261_r;
      node1266_r = node1260_r & pixel[287];
      node1266_l = node1260_r & ~pixel[287];
      node1267_r = node1266_l & pixel[149];
      node1267_l = node1266_l & ~pixel[149];
      node1268 = node1267_l;
      node1269 = node1267_r;
      node1270_r = node1266_r & pixel[326];
      node1270_l = node1266_r & ~pixel[326];
      node1271 = node1270_l;
      node1272 = node1270_r;
      node1273_r = node1259_r & pixel[209];
      node1273_l = node1259_r & ~pixel[209];
      node1274_r = node1273_l & pixel[206];
      node1274_l = node1273_l & ~pixel[206];
      node1275 = node1274_l;
      node1276_r = node1274_r & pixel[159];
      node1276_l = node1274_r & ~pixel[159];
      node1277 = node1276_l;
      node1278 = node1276_r;
      node1279_r = node1273_r & pixel[271];
      node1279_l = node1273_r & ~pixel[271];
      node1280_r = node1279_l & pixel[270];
      node1280_l = node1279_l & ~pixel[270];
      node1281 = node1280_l;
      node1282 = node1280_r;
      node1283_r = node1279_r & pixel[349];
      node1283_l = node1279_r & ~pixel[349];
      node1284 = node1283_l;
      node1285 = node1283_r;
      node1286_r = node1258_r & pixel[484];
      node1286_l = node1258_r & ~pixel[484];
      node1287_r = node1286_l & pixel[158];
      node1287_l = node1286_l & ~pixel[158];
      node1288_r = node1287_l & pixel[580];
      node1288_l = node1287_l & ~pixel[580];
      node1289_r = node1288_l & pixel[181];
      node1289_l = node1288_l & ~pixel[181];
      node1290 = node1289_l;
      node1291 = node1289_r;
      node1292_r = node1288_r & pixel[270];
      node1292_l = node1288_r & ~pixel[270];
      node1293 = node1292_l;
      node1294 = node1292_r;
      node1295_r = node1287_r & pixel[299];
      node1295_l = node1287_r & ~pixel[299];
      node1296_r = node1295_l & pixel[294];
      node1296_l = node1295_l & ~pixel[294];
      node1297 = node1296_l;
      node1298 = node1296_r;
      node1299_r = node1295_r & pixel[324];
      node1299_l = node1295_r & ~pixel[324];
      node1300 = node1299_l;
      node1301 = node1299_r;
      node1302_r = node1286_r & pixel[379];
      node1302_l = node1286_r & ~pixel[379];
      node1303_r = node1302_l & pixel[299];
      node1303_l = node1302_l & ~pixel[299];
      node1304_r = node1303_l & pixel[657];
      node1304_l = node1303_l & ~pixel[657];
      node1305 = node1304_l;
      node1306 = node1304_r;
      node1307_r = node1303_r & pixel[175];
      node1307_l = node1303_r & ~pixel[175];
      node1308 = node1307_l;
      node1309 = node1307_r;
      node1310_r = node1302_r & pixel[485];
      node1310_l = node1302_r & ~pixel[485];
      node1311_r = node1310_l & pixel[272];
      node1311_l = node1310_l & ~pixel[272];
      node1312 = node1311_l;
      node1313 = node1311_r;
      node1314_r = node1310_r & pixel[543];
      node1314_l = node1310_r & ~pixel[543];
      node1315 = node1314_l;
      node1316 = node1314_r;
      node1317_r = node1257_r & pixel[629];
      node1317_l = node1257_r & ~pixel[629];
      node1318_r = node1317_l & pixel[470];
      node1318_l = node1317_l & ~pixel[470];
      node1319_r = node1318_l & pixel[213];
      node1319_l = node1318_l & ~pixel[213];
      node1320_r = node1319_l & pixel[379];
      node1320_l = node1319_l & ~pixel[379];
      node1321 = node1320_l;
      node1322_r = node1320_r & pixel[542];
      node1322_l = node1320_r & ~pixel[542];
      node1323 = node1322_l;
      node1324 = node1322_r;
      node1325_r = node1319_r & pixel[428];
      node1325_l = node1319_r & ~pixel[428];
      node1326_r = node1325_l & pixel[150];
      node1326_l = node1325_l & ~pixel[150];
      node1327 = node1326_l;
      node1328 = node1326_r;
      node1329_r = node1325_r & pixel[511];
      node1329_l = node1325_r & ~pixel[511];
      node1330 = node1329_l;
      node1331 = node1329_r;
      node1332_r = node1318_r & pixel[271];
      node1332_l = node1318_r & ~pixel[271];
      node1333_r = node1332_l & pixel[269];
      node1333_l = node1332_l & ~pixel[269];
      node1334_r = node1333_l & pixel[541];
      node1334_l = node1333_l & ~pixel[541];
      node1335 = node1334_l;
      node1336 = node1334_r;
      node1337 = node1333_r;
      node1338_r = node1332_r & pixel[406];
      node1338_l = node1332_r & ~pixel[406];
      node1339 = node1338_l;
      node1340_r = node1338_r & pixel[444];
      node1340_l = node1338_r & ~pixel[444];
      node1341 = node1340_l;
      node1342 = node1340_r;
      node1343_r = node1317_r & pixel[244];
      node1343_l = node1317_r & ~pixel[244];
      node1344_r = node1343_l & pixel[463];
      node1344_l = node1343_l & ~pixel[463];
      node1345_r = node1344_l & pixel[298];
      node1345_l = node1344_l & ~pixel[298];
      node1346_r = node1345_l & pixel[662];
      node1346_l = node1345_l & ~pixel[662];
      node1347 = node1346_l;
      node1348 = node1346_r;
      node1349_r = node1345_r & pixel[378];
      node1349_l = node1345_r & ~pixel[378];
      node1350 = node1349_l;
      node1351 = node1349_r;
      node1352_r = node1344_r & pixel[412];
      node1352_l = node1344_r & ~pixel[412];
      node1353_r = node1352_l & pixel[386];
      node1353_l = node1352_l & ~pixel[386];
      node1354 = node1353_l;
      node1355 = node1353_r;
      node1356_r = node1352_r & pixel[268];
      node1356_l = node1352_r & ~pixel[268];
      node1357 = node1356_l;
      node1358 = node1356_r;
      node1359_r = node1343_r & pixel[661];
      node1359_l = node1343_r & ~pixel[661];
      node1360_r = node1359_l & pixel[625];
      node1360_l = node1359_l & ~pixel[625];
      node1361_r = node1360_l & pixel[186];
      node1361_l = node1360_l & ~pixel[186];
      node1362 = node1361_l;
      node1363 = node1361_r;
      node1364_r = node1360_r & pixel[408];
      node1364_l = node1360_r & ~pixel[408];
      node1365 = node1364_l;
      node1366 = node1364_r;
      node1367_r = node1359_r & pixel[404];
      node1367_l = node1359_r & ~pixel[404];
      node1368_r = node1367_l & pixel[541];
      node1368_l = node1367_l & ~pixel[541];
      node1369 = node1368_l;
      node1370 = node1368_r;
      node1371_r = node1367_r & pixel[355];
      node1371_l = node1367_r & ~pixel[355];
      node1372 = node1371_l;
      node1373 = node1371_r;
      node1374_r = node910_r & pixel[686];
      node1374_l = node910_r & ~pixel[686];
      node1375_r = node1374_l & pixel[322];
      node1375_l = node1374_l & ~pixel[322];
      node1376_r = node1375_l & pixel[215];
      node1376_l = node1375_l & ~pixel[215];
      node1377_r = node1376_l & pixel[213];
      node1377_l = node1376_l & ~pixel[213];
      node1378_r = node1377_l & pixel[656];
      node1378_l = node1377_l & ~pixel[656];
      node1379_r = node1378_l & pixel[537];
      node1379_l = node1378_l & ~pixel[537];
      node1380_r = node1379_l & pixel[268];
      node1380_l = node1379_l & ~pixel[268];
      node1381_r = node1380_l & pixel[660];
      node1381_l = node1380_l & ~pixel[660];
      node1382 = node1381_l;
      node1383 = node1381_r;
      node1384_r = node1380_r & pixel[123];
      node1384_l = node1380_r & ~pixel[123];
      node1385 = node1384_l;
      node1386 = node1384_r;
      node1387_r = node1379_r & pixel[496];
      node1387_l = node1379_r & ~pixel[496];
      node1388_r = node1387_l & pixel[320];
      node1388_l = node1387_l & ~pixel[320];
      node1389 = node1388_l;
      node1390 = node1388_r;
      node1391_r = node1387_r & pixel[162];
      node1391_l = node1387_r & ~pixel[162];
      node1392 = node1391_l;
      node1393 = node1391_r;
      node1394_r = node1378_r & pixel[327];
      node1394_l = node1378_r & ~pixel[327];
      node1395_r = node1394_l & pixel[268];
      node1395_l = node1394_l & ~pixel[268];
      node1396_r = node1395_l & pixel[658];
      node1396_l = node1395_l & ~pixel[658];
      node1397 = node1396_l;
      node1398 = node1396_r;
      node1399_r = node1395_r & pixel[237];
      node1399_l = node1395_r & ~pixel[237];
      node1400 = node1399_l;
      node1401 = node1399_r;
      node1402_r = node1394_r & pixel[378];
      node1402_l = node1394_r & ~pixel[378];
      node1403_r = node1402_l & pixel[603];
      node1403_l = node1402_l & ~pixel[603];
      node1404 = node1403_l;
      node1405 = node1403_r;
      node1406_r = node1402_r & pixel[157];
      node1406_l = node1402_r & ~pixel[157];
      node1407 = node1406_l;
      node1408 = node1406_r;
      node1409_r = node1377_r & pixel[296];
      node1409_l = node1377_r & ~pixel[296];
      node1410_r = node1409_l & pixel[319];
      node1410_l = node1409_l & ~pixel[319];
      node1411_r = node1410_l & pixel[402];
      node1411_l = node1410_l & ~pixel[402];
      node1412_r = node1411_l & pixel[344];
      node1412_l = node1411_l & ~pixel[344];
      node1413 = node1412_l;
      node1414 = node1412_r;
      node1415_r = node1411_r & pixel[316];
      node1415_l = node1411_r & ~pixel[316];
      node1416 = node1415_l;
      node1417 = node1415_r;
      node1418_r = node1410_r & pixel[524];
      node1418_l = node1410_r & ~pixel[524];
      node1419_r = node1418_l & pixel[495];
      node1419_l = node1418_l & ~pixel[495];
      node1420 = node1419_l;
      node1421 = node1419_r;
      node1422_r = node1418_r & pixel[321];
      node1422_l = node1418_r & ~pixel[321];
      node1423 = node1422_l;
      node1424 = node1422_r;
      node1425_r = node1409_r & pixel[661];
      node1425_l = node1409_r & ~pixel[661];
      node1426_r = node1425_l & pixel[344];
      node1426_l = node1425_l & ~pixel[344];
      node1427_r = node1426_l & pixel[321];
      node1427_l = node1426_l & ~pixel[321];
      node1428 = node1427_l;
      node1429 = node1427_r;
      node1430_r = node1426_r & pixel[399];
      node1430_l = node1426_r & ~pixel[399];
      node1431 = node1430_l;
      node1432 = node1430_r;
      node1433_r = node1425_r & pixel[125];
      node1433_l = node1425_r & ~pixel[125];
      node1434_r = node1433_l & pixel[153];
      node1434_l = node1433_l & ~pixel[153];
      node1435 = node1434_l;
      node1436 = node1434_r;
      node1437_r = node1433_r & pixel[404];
      node1437_l = node1433_r & ~pixel[404];
      node1438 = node1437_l;
      node1439 = node1437_r;
      node1440_r = node1376_r & pixel[346];
      node1440_l = node1376_r & ~pixel[346];
      node1441_r = node1440_l & pixel[320];
      node1441_l = node1440_l & ~pixel[320];
      node1442_r = node1441_l & pixel[126];
      node1442_l = node1441_l & ~pixel[126];
      node1443_r = node1442_l & pixel[315];
      node1443_l = node1442_l & ~pixel[315];
      node1444_r = node1443_l & pixel[653];
      node1444_l = node1443_l & ~pixel[653];
      node1445 = node1444_l;
      node1446 = node1444_r;
      node1447_r = node1443_r & pixel[402];
      node1447_l = node1443_r & ~pixel[402];
      node1448 = node1447_l;
      node1449 = node1447_r;
      node1450_r = node1442_r & pixel[374];
      node1450_l = node1442_r & ~pixel[374];
      node1451_r = node1450_l & pixel[369];
      node1451_l = node1450_l & ~pixel[369];
      node1452 = node1451_l;
      node1453 = node1451_r;
      node1454_r = node1450_r & pixel[544];
      node1454_l = node1450_r & ~pixel[544];
      node1455 = node1454_l;
      node1456 = node1454_r;
      node1457_r = node1441_r & pixel[348];
      node1457_l = node1441_r & ~pixel[348];
      node1458_r = node1457_l & pixel[656];
      node1458_l = node1457_l & ~pixel[656];
      node1459 = node1458_l;
      node1460_r = node1458_r & pixel[681];
      node1460_l = node1458_r & ~pixel[681];
      node1461 = node1460_l;
      node1462 = node1460_r;
      node1463_r = node1457_r & pixel[406];
      node1463_l = node1457_r & ~pixel[406];
      node1464_r = node1463_l & pixel[595];
      node1464_l = node1463_l & ~pixel[595];
      node1465 = node1464_l;
      node1466 = node1464_r;
      node1467_r = node1463_r & pixel[465];
      node1467_l = node1463_r & ~pixel[465];
      node1468 = node1467_l;
      node1469 = node1467_r;
      node1470_r = node1440_r & pixel[457];
      node1470_l = node1440_r & ~pixel[457];
      node1471_r = node1470_l & pixel[371];
      node1471_l = node1470_l & ~pixel[371];
      node1472_r = node1471_l & pixel[375];
      node1472_l = node1471_l & ~pixel[375];
      node1473_r = node1472_l & pixel[546];
      node1473_l = node1472_l & ~pixel[546];
      node1474 = node1473_l;
      node1475 = node1473_r;
      node1476_r = node1472_r & pixel[299];
      node1476_l = node1472_r & ~pixel[299];
      node1477 = node1476_l;
      node1478 = node1476_r;
      node1479_r = node1471_r & pixel[260];
      node1479_l = node1471_r & ~pixel[260];
      node1480_r = node1479_l & pixel[330];
      node1480_l = node1479_l & ~pixel[330];
      node1481 = node1480_l;
      node1482 = node1480_r;
      node1483_r = node1479_r & pixel[464];
      node1483_l = node1479_r & ~pixel[464];
      node1484 = node1483_l;
      node1485 = node1483_r;
      node1486_r = node1470_r & pixel[495];
      node1486_l = node1470_r & ~pixel[495];
      node1487_r = node1486_l & pixel[378];
      node1487_l = node1486_l & ~pixel[378];
      node1488_r = node1487_l & pixel[129];
      node1488_l = node1487_l & ~pixel[129];
      node1489 = node1488_l;
      node1490 = node1488_r;
      node1491_r = node1487_r & pixel[372];
      node1491_l = node1487_r & ~pixel[372];
      node1492 = node1491_l;
      node1493 = node1491_r;
      node1494_r = node1486_r & pixel[603];
      node1494_l = node1486_r & ~pixel[603];
      node1495_r = node1494_l & pixel[597];
      node1495_l = node1494_l & ~pixel[597];
      node1496 = node1495_l;
      node1497 = node1495_r;
      node1498_r = node1494_r & pixel[102];
      node1498_l = node1494_r & ~pixel[102];
      node1499 = node1498_l;
      node1500 = node1498_r;
      node1501_r = node1375_r & pixel[402];
      node1501_l = node1375_r & ~pixel[402];
      node1502_r = node1501_l & pixel[180];
      node1502_l = node1501_l & ~pixel[180];
      node1503_r = node1502_l & pixel[267];
      node1503_l = node1502_l & ~pixel[267];
      node1504_r = node1503_l & pixel[514];
      node1504_l = node1503_l & ~pixel[514];
      node1505_r = node1504_l & pixel[160];
      node1505_l = node1504_l & ~pixel[160];
      node1506_r = node1505_l & pixel[435];
      node1506_l = node1505_l & ~pixel[435];
      node1507 = node1506_l;
      node1508 = node1506_r;
      node1509 = node1505_r;
      node1510_r = node1504_r & pixel[466];
      node1510_l = node1504_r & ~pixel[466];
      node1511_r = node1510_l & pixel[553];
      node1511_l = node1510_l & ~pixel[553];
      node1512 = node1511_l;
      node1513 = node1511_r;
      node1514_r = node1510_r & pixel[270];
      node1514_l = node1510_r & ~pixel[270];
      node1515 = node1514_l;
      node1516 = node1514_r;
      node1517_r = node1503_r & pixel[409];
      node1517_l = node1503_r & ~pixel[409];
      node1518_r = node1517_l & pixel[580];
      node1518_l = node1517_l & ~pixel[580];
      node1519_r = node1518_l & pixel[550];
      node1519_l = node1518_l & ~pixel[550];
      node1520 = node1519_l;
      node1521 = node1519_r;
      node1522_r = node1518_r & pixel[101];
      node1522_l = node1518_r & ~pixel[101];
      node1523 = node1522_l;
      node1524 = node1522_r;
      node1525_r = node1517_r & pixel[512];
      node1525_l = node1517_r & ~pixel[512];
      node1526_r = node1525_l & pixel[550];
      node1526_l = node1525_l & ~pixel[550];
      node1527 = node1526_l;
      node1528 = node1526_r;
      node1529_r = node1525_r & pixel[654];
      node1529_l = node1525_r & ~pixel[654];
      node1530 = node1529_l;
      node1531 = node1529_r;
      node1532_r = node1502_r & pixel[326];
      node1532_l = node1502_r & ~pixel[326];
      node1533_r = node1532_l & pixel[542];
      node1533_l = node1532_l & ~pixel[542];
      node1534_r = node1533_l & pixel[550];
      node1534_l = node1533_l & ~pixel[550];
      node1535_r = node1534_l & pixel[241];
      node1535_l = node1534_l & ~pixel[241];
      node1536 = node1535_l;
      node1537 = node1535_r;
      node1538_r = node1534_r & pixel[538];
      node1538_l = node1534_r & ~pixel[538];
      node1539 = node1538_l;
      node1540 = node1538_r;
      node1541_r = node1533_r & pixel[240];
      node1541_l = node1533_r & ~pixel[240];
      node1542_r = node1541_l & pixel[316];
      node1542_l = node1541_l & ~pixel[316];
      node1543 = node1542_l;
      node1544 = node1542_r;
      node1545_r = node1541_r & pixel[292];
      node1545_l = node1541_r & ~pixel[292];
      node1546 = node1545_l;
      node1547 = node1545_r;
      node1548_r = node1532_r & pixel[348];
      node1548_l = node1532_r & ~pixel[348];
      node1549_r = node1548_l & pixel[635];
      node1549_l = node1548_l & ~pixel[635];
      node1550_r = node1549_l & pixel[514];
      node1550_l = node1549_l & ~pixel[514];
      node1551 = node1550_l;
      node1552 = node1550_r;
      node1553_r = node1549_r & pixel[412];
      node1553_l = node1549_r & ~pixel[412];
      node1554 = node1553_l;
      node1555 = node1553_r;
      node1556_r = node1548_r & pixel[433];
      node1556_l = node1548_r & ~pixel[433];
      node1557_r = node1556_l & pixel[240];
      node1557_l = node1556_l & ~pixel[240];
      node1558 = node1557_l;
      node1559 = node1557_r;
      node1560_r = node1556_r & pixel[526];
      node1560_l = node1556_r & ~pixel[526];
      node1561 = node1560_l;
      node1562 = node1560_r;
      node1563_r = node1501_r & pixel[296];
      node1563_l = node1501_r & ~pixel[296];
      node1564_r = node1563_l & pixel[494];
      node1564_l = node1563_l & ~pixel[494];
      node1565_r = node1564_l & pixel[271];
      node1565_l = node1564_l & ~pixel[271];
      node1566_r = node1565_l & pixel[544];
      node1566_l = node1565_l & ~pixel[544];
      node1567_r = node1566_l & pixel[384];
      node1567_l = node1566_l & ~pixel[384];
      node1568 = node1567_l;
      node1569 = node1567_r;
      node1570_r = node1566_r & pixel[260];
      node1570_l = node1566_r & ~pixel[260];
      node1571 = node1570_l;
      node1572 = node1570_r;
      node1573_r = node1565_r & pixel[630];
      node1573_l = node1565_r & ~pixel[630];
      node1574_r = node1573_l & pixel[378];
      node1574_l = node1573_l & ~pixel[378];
      node1575 = node1574_l;
      node1576 = node1574_r;
      node1577_r = node1573_r & pixel[538];
      node1577_l = node1573_r & ~pixel[538];
      node1578 = node1577_l;
      node1579 = node1577_r;
      node1580_r = node1564_r & pixel[130];
      node1580_l = node1564_r & ~pixel[130];
      node1581_r = node1580_l & pixel[99];
      node1581_l = node1580_l & ~pixel[99];
      node1582_r = node1581_l & pixel[186];
      node1582_l = node1581_l & ~pixel[186];
      node1583 = node1582_l;
      node1584 = node1582_r;
      node1585_r = node1581_r & pixel[594];
      node1585_l = node1581_r & ~pixel[594];
      node1586 = node1585_l;
      node1587 = node1585_r;
      node1588_r = node1580_r & pixel[648];
      node1588_l = node1580_r & ~pixel[648];
      node1589_r = node1588_l & pixel[273];
      node1589_l = node1588_l & ~pixel[273];
      node1590 = node1589_l;
      node1591 = node1589_r;
      node1592 = node1588_r;
      node1593_r = node1563_r & pixel[659];
      node1593_l = node1563_r & ~pixel[659];
      node1594_r = node1593_l & pixel[528];
      node1594_l = node1593_l & ~pixel[528];
      node1595_r = node1594_l & pixel[654];
      node1595_l = node1594_l & ~pixel[654];
      node1596_r = node1595_l & pixel[383];
      node1596_l = node1595_l & ~pixel[383];
      node1597 = node1596_l;
      node1598 = node1596_r;
      node1599_r = node1595_r & pixel[293];
      node1599_l = node1595_r & ~pixel[293];
      node1600 = node1599_l;
      node1601 = node1599_r;
      node1602_r = node1594_r & pixel[385];
      node1602_l = node1594_r & ~pixel[385];
      node1603_r = node1602_l & pixel[553];
      node1603_l = node1602_l & ~pixel[553];
      node1604 = node1603_l;
      node1605 = node1603_r;
      node1606_r = node1602_r & pixel[387];
      node1606_l = node1602_r & ~pixel[387];
      node1607 = node1606_l;
      node1608 = node1606_r;
      node1609_r = node1593_r & pixel[656];
      node1609_l = node1593_r & ~pixel[656];
      node1610_r = node1609_l & pixel[581];
      node1610_l = node1609_l & ~pixel[581];
      node1611_r = node1610_l & pixel[458];
      node1611_l = node1610_l & ~pixel[458];
      node1612 = node1611_l;
      node1613 = node1611_r;
      node1614_r = node1610_r & pixel[401];
      node1614_l = node1610_r & ~pixel[401];
      node1615 = node1614_l;
      node1616 = node1614_r;
      node1617_r = node1609_r & pixel[610];
      node1617_l = node1609_r & ~pixel[610];
      node1618_r = node1617_l & pixel[485];
      node1618_l = node1617_l & ~pixel[485];
      node1619 = node1618_l;
      node1620 = node1618_r;
      node1621_r = node1617_r & pixel[466];
      node1621_l = node1617_r & ~pixel[466];
      node1622 = node1621_l;
      node1623 = node1621_r;
      node1624_r = node1374_r & pixel[262];
      node1624_l = node1374_r & ~pixel[262];
      node1625_r = node1624_l & pixel[403];
      node1625_l = node1624_l & ~pixel[403];
      node1626_r = node1625_l & pixel[486];
      node1626_l = node1625_l & ~pixel[486];
      node1627_r = node1626_l & pixel[267];
      node1627_l = node1626_l & ~pixel[267];
      node1628_r = node1627_l & pixel[149];
      node1628_l = node1627_l & ~pixel[149];
      node1629_r = node1628_l & pixel[595];
      node1629_l = node1628_l & ~pixel[595];
      node1630_r = node1629_l & pixel[571];
      node1630_l = node1629_l & ~pixel[571];
      node1631 = node1630_l;
      node1632 = node1630_r;
      node1633 = node1629_r;
      node1634_r = node1628_r & pixel[209];
      node1634_l = node1628_r & ~pixel[209];
      node1635_r = node1634_l & pixel[546];
      node1635_l = node1634_l & ~pixel[546];
      node1636 = node1635_l;
      node1637 = node1635_r;
      node1638_r = node1634_r & pixel[575];
      node1638_l = node1634_r & ~pixel[575];
      node1639 = node1638_l;
      node1640 = node1638_r;
      node1641_r = node1627_r & pixel[608];
      node1641_l = node1627_r & ~pixel[608];
      node1642_r = node1641_l & pixel[294];
      node1642_l = node1641_l & ~pixel[294];
      node1643_r = node1642_l & pixel[297];
      node1643_l = node1642_l & ~pixel[297];
      node1644 = node1643_l;
      node1645 = node1643_r;
      node1646_r = node1642_r & pixel[551];
      node1646_l = node1642_r & ~pixel[551];
      node1647 = node1646_l;
      node1648 = node1646_r;
      node1649_r = node1641_r & pixel[605];
      node1649_l = node1641_r & ~pixel[605];
      node1650 = node1649_l;
      node1651_r = node1649_r & pixel[600];
      node1651_l = node1649_r & ~pixel[600];
      node1652 = node1651_l;
      node1653 = node1651_r;
      node1654_r = node1626_r & pixel[662];
      node1654_l = node1626_r & ~pixel[662];
      node1655_r = node1654_l & pixel[466];
      node1655_l = node1654_l & ~pixel[466];
      node1656_r = node1655_l & pixel[346];
      node1656_l = node1655_l & ~pixel[346];
      node1657_r = node1656_l & pixel[237];
      node1657_l = node1656_l & ~pixel[237];
      node1658 = node1657_l;
      node1659 = node1657_r;
      node1660_r = node1656_r & pixel[568];
      node1660_l = node1656_r & ~pixel[568];
      node1661 = node1660_l;
      node1662 = node1660_r;
      node1663_r = node1655_r & pixel[207];
      node1663_l = node1655_r & ~pixel[207];
      node1664_r = node1663_l & pixel[682];
      node1664_l = node1663_l & ~pixel[682];
      node1665 = node1664_l;
      node1666 = node1664_r;
      node1667_r = node1663_r & pixel[483];
      node1667_l = node1663_r & ~pixel[483];
      node1668 = node1667_l;
      node1669 = node1667_r;
      node1670_r = node1654_r & pixel[538];
      node1670_l = node1654_r & ~pixel[538];
      node1671_r = node1670_l & pixel[345];
      node1671_l = node1670_l & ~pixel[345];
      node1672_r = node1671_l & pixel[498];
      node1672_l = node1671_l & ~pixel[498];
      node1673 = node1672_l;
      node1674 = node1672_r;
      node1675_r = node1671_r & pixel[527];
      node1675_l = node1671_r & ~pixel[527];
      node1676 = node1675_l;
      node1677 = node1675_r;
      node1678_r = node1670_r & pixel[585];
      node1678_l = node1670_r & ~pixel[585];
      node1679 = node1678_l;
      node1680 = node1678_r;
      node1681_r = node1625_r & pixel[350];
      node1681_l = node1625_r & ~pixel[350];
      node1682_r = node1681_l & pixel[599];
      node1682_l = node1681_l & ~pixel[599];
      node1683_r = node1682_l & pixel[514];
      node1683_l = node1682_l & ~pixel[514];
      node1684_r = node1683_l & pixel[215];
      node1684_l = node1683_l & ~pixel[215];
      node1685_r = node1684_l & pixel[681];
      node1685_l = node1684_l & ~pixel[681];
      node1686 = node1685_l;
      node1687 = node1685_r;
      node1688_r = node1684_r & pixel[553];
      node1688_l = node1684_r & ~pixel[553];
      node1689 = node1688_l;
      node1690 = node1688_r;
      node1691_r = node1683_r & pixel[329];
      node1691_l = node1683_r & ~pixel[329];
      node1692_r = node1691_l & pixel[457];
      node1692_l = node1691_l & ~pixel[457];
      node1693 = node1692_l;
      node1694 = node1692_r;
      node1695 = node1691_r;
      node1696_r = node1682_r & pixel[293];
      node1696_l = node1682_r & ~pixel[293];
      node1697_r = node1696_l & pixel[470];
      node1697_l = node1696_l & ~pixel[470];
      node1698_r = node1697_l & pixel[515];
      node1698_l = node1697_l & ~pixel[515];
      node1699 = node1698_l;
      node1700 = node1698_r;
      node1701_r = node1697_r & pixel[313];
      node1701_l = node1697_r & ~pixel[313];
      node1702 = node1701_l;
      node1703 = node1701_r;
      node1704_r = node1696_r & pixel[406];
      node1704_l = node1696_r & ~pixel[406];
      node1705_r = node1704_l & pixel[328];
      node1705_l = node1704_l & ~pixel[328];
      node1706 = node1705_l;
      node1707 = node1705_r;
      node1708_r = node1704_r & pixel[683];
      node1708_l = node1704_r & ~pixel[683];
      node1709 = node1708_l;
      node1710 = node1708_r;
      node1711_r = node1681_r & pixel[326];
      node1711_l = node1681_r & ~pixel[326];
      node1712_r = node1711_l & pixel[345];
      node1712_l = node1711_l & ~pixel[345];
      node1713_r = node1712_l & pixel[522];
      node1713_l = node1712_l & ~pixel[522];
      node1714_r = node1713_l & pixel[293];
      node1714_l = node1713_l & ~pixel[293];
      node1715 = node1714_l;
      node1716 = node1714_r;
      node1717_r = node1713_r & pixel[551];
      node1717_l = node1713_r & ~pixel[551];
      node1718 = node1717_l;
      node1719 = node1717_r;
      node1720_r = node1712_r & pixel[208];
      node1720_l = node1712_r & ~pixel[208];
      node1721_r = node1720_l & pixel[689];
      node1721_l = node1720_l & ~pixel[689];
      node1722 = node1721_l;
      node1723 = node1721_r;
      node1724_r = node1720_r & pixel[172];
      node1724_l = node1720_r & ~pixel[172];
      node1725 = node1724_l;
      node1726 = node1724_r;
      node1727_r = node1711_r & pixel[177];
      node1727_l = node1711_r & ~pixel[177];
      node1728_r = node1727_l & pixel[494];
      node1728_l = node1727_l & ~pixel[494];
      node1729 = node1728_l;
      node1730_r = node1728_r & pixel[573];
      node1730_l = node1728_r & ~pixel[573];
      node1731 = node1730_l;
      node1732 = node1730_r;
      node1733_r = node1727_r & pixel[689];
      node1733_l = node1727_r & ~pixel[689];
      node1734_r = node1733_l & pixel[346];
      node1734_l = node1733_l & ~pixel[346];
      node1735 = node1734_l;
      node1736 = node1734_r;
      node1737_r = node1733_r & pixel[543];
      node1737_l = node1733_r & ~pixel[543];
      node1738 = node1737_l;
      node1739 = node1737_r;
      node1740_r = node1624_r & pixel[456];
      node1740_l = node1624_r & ~pixel[456];
      node1741_r = node1740_l & pixel[407];
      node1741_l = node1740_l & ~pixel[407];
      node1742_r = node1741_l & pixel[190];
      node1742_l = node1741_l & ~pixel[190];
      node1743_r = node1742_l & pixel[513];
      node1743_l = node1742_l & ~pixel[513];
      node1744_r = node1743_l & pixel[355];
      node1744_l = node1743_l & ~pixel[355];
      node1745_r = node1744_l & pixel[323];
      node1745_l = node1744_l & ~pixel[323];
      node1746 = node1745_l;
      node1747 = node1745_r;
      node1748_r = node1744_r & pixel[158];
      node1748_l = node1744_r & ~pixel[158];
      node1749 = node1748_l;
      node1750 = node1748_r;
      node1751_r = node1743_r & pixel[440];
      node1751_l = node1743_r & ~pixel[440];
      node1752_r = node1751_l & pixel[158];
      node1752_l = node1751_l & ~pixel[158];
      node1753 = node1752_l;
      node1754 = node1752_r;
      node1755_r = node1751_r & pixel[425];
      node1755_l = node1751_r & ~pixel[425];
      node1756 = node1755_l;
      node1757 = node1755_r;
      node1758_r = node1742_r & pixel[297];
      node1758_l = node1742_r & ~pixel[297];
      node1759_r = node1758_l & pixel[328];
      node1759_l = node1758_l & ~pixel[328];
      node1760 = node1759_l;
      node1761 = node1759_r;
      node1762_r = node1758_r & pixel[322];
      node1762_l = node1758_r & ~pixel[322];
      node1763 = node1762_l;
      node1764 = node1762_r;
      node1765_r = node1741_r & pixel[537];
      node1765_l = node1741_r & ~pixel[537];
      node1766_r = node1765_l & pixel[611];
      node1766_l = node1765_l & ~pixel[611];
      node1767_r = node1766_l & pixel[433];
      node1767_l = node1766_l & ~pixel[433];
      node1768_r = node1767_l & pixel[323];
      node1768_l = node1767_l & ~pixel[323];
      node1769 = node1768_l;
      node1770 = node1768_r;
      node1771_r = node1767_r & pixel[380];
      node1771_l = node1767_r & ~pixel[380];
      node1772 = node1771_l;
      node1773 = node1771_r;
      node1774_r = node1766_r & pixel[468];
      node1774_l = node1766_r & ~pixel[468];
      node1775_r = node1774_l & pixel[373];
      node1775_l = node1774_l & ~pixel[373];
      node1776 = node1775_l;
      node1777 = node1775_r;
      node1778 = node1774_r;
      node1779_r = node1765_r & pixel[162];
      node1779_l = node1765_r & ~pixel[162];
      node1780 = node1779_l;
      node1781 = node1779_r;
      node1782_r = node1740_r & pixel[273];
      node1782_l = node1740_r & ~pixel[273];
      node1783_r = node1782_l & pixel[290];
      node1783_l = node1782_l & ~pixel[290];
      node1784_r = node1783_l & pixel[542];
      node1784_l = node1783_l & ~pixel[542];
      node1785 = node1784_l;
      node1786_r = node1784_r & pixel[371];
      node1786_l = node1784_r & ~pixel[371];
      node1787 = node1786_l;
      node1788 = node1786_r;
      node1789_r = node1783_r & pixel[581];
      node1789_l = node1783_r & ~pixel[581];
      node1790_r = node1789_l & pixel[326];
      node1790_l = node1789_l & ~pixel[326];
      node1791_r = node1790_l & pixel[157];
      node1791_l = node1790_l & ~pixel[157];
      node1792 = node1791_l;
      node1793 = node1791_r;
      node1794_r = node1790_r & pixel[322];
      node1794_l = node1790_r & ~pixel[322];
      node1795 = node1794_l;
      node1796 = node1794_r;
      node1797_r = node1789_r & pixel[324];
      node1797_l = node1789_r & ~pixel[324];
      node1798_r = node1797_l & pixel[662];
      node1798_l = node1797_l & ~pixel[662];
      node1799 = node1798_l;
      node1800 = node1798_r;
      node1801_r = node1797_r & pixel[319];
      node1801_l = node1797_r & ~pixel[319];
      node1802 = node1801_l;
      node1803 = node1801_r;
      node1804_r = node1782_r & pixel[442];
      node1804_l = node1782_r & ~pixel[442];
      node1805_r = node1804_l & pixel[627];
      node1805_l = node1804_l & ~pixel[627];
      node1806_r = node1805_l & pixel[292];
      node1806_l = node1805_l & ~pixel[292];
      node1807_r = node1806_l & pixel[288];
      node1807_l = node1806_l & ~pixel[288];
      node1808 = node1807_l;
      node1809 = node1807_r;
      node1810_r = node1806_r & pixel[157];
      node1810_l = node1806_r & ~pixel[157];
      node1811 = node1810_l;
      node1812 = node1810_r;
      node1813_r = node1805_r & pixel[379];
      node1813_l = node1805_r & ~pixel[379];
      node1814_r = node1813_l & pixel[436];
      node1814_l = node1813_l & ~pixel[436];
      node1815 = node1814_l;
      node1816 = node1814_r;
      node1817_r = node1813_r & pixel[347];
      node1817_l = node1813_r & ~pixel[347];
      node1818 = node1817_l;
      node1819 = node1817_r;
      node1820_r = node1804_r & pixel[498];
      node1820_l = node1804_r & ~pixel[498];
      node1821_r = node1820_l & pixel[436];
      node1821_l = node1820_l & ~pixel[436];
      node1822 = node1821_l;
      node1823_r = node1821_r & pixel[345];
      node1823_l = node1821_r & ~pixel[345];
      node1824 = node1823_l;
      node1825 = node1823_r;
      node1826_r = node1820_r & pixel[369];
      node1826_l = node1820_r & ~pixel[369];
      node1827_r = node1826_l & pixel[489];
      node1827_l = node1826_l & ~pixel[489];
      node1828 = node1827_l;
      node1829 = node1827_r;
      node1830 = node1826_r;
      result0 = node21 | node29 | node42 | node45 | node70 | node78 | node113 | node153 | node157 | node168 | node182 | node192 | node200 | node206 | node211 | node217 | node232 | node236 | node273 | node278 | node288 | node303 | node307 | node339 | node378 | node419 | node424 | node430 | node432 | node437 | node446 | node496 | node501 | node515 | node521 | node522 | node537 | node538 | node544 | node559 | node592 | node633 | node651 | node752 | node772 | node774 | node775 | node790 | node805 | node832 | node860 | node875 | node883 | node887 | node890 | node894 | node908 | node909 | node927 | node935 | node965 | node969 | node1007 | node1022 | node1023 | node1025 | node1034 | node1041 | node1064 | node1065 | node1069 | node1093 | node1142 | node1173 | node1174 | node1189 | node1191 | node1196 | node1200 | node1207 | node1211 | node1214 | node1215 | node1217 | node1218 | node1229 | node1234 | node1236 | node1241 | node1252 | node1253 | node1282 | node1284 | node1308 | node1339 | node1350 | node1365 | node1366 | node1369 | node1370 | node1482 | node1499 | node1591 | node1601 | node1707 | node1756 | node1796 | node1815 | node1822 | node1825 | node1828;
      result1 = node13 | node35 | node48 | node49 | node62 | node225 | node226 | node243 | node380 | node406 | node409 | node414 | node418 | node566 | node570 | node919 | node920 | node929 | node938 | node977 | node992 | node1097 | node1162 | node1507 | node1520 | node1527 | node1536 | node1537 | node1644 | node1647 | node1666 | node1716;
      result2 = node25 | node41 | node56 | node63 | node69 | node75 | node83 | node89 | node137 | node139 | node181 | node184 | node203 | node213 | node216 | node235 | node247 | node255 | node261 | node262 | node265 | node305 | node354 | node365 | node368 | node384 | node387 | node404 | node445 | node477 | node486 | node543 | node551 | node629 | node636 | node637 | node677 | node768 | node784 | node821 | node828 | node837 | node840 | node856 | node886 | node893 | node899 | node941 | node943 | node958 | node959 | node963 | node964 | node968 | node980 | node1008 | node1035 | node1038 | node1040 | node1048 | node1049 | node1062 | node1068 | node1071 | node1072 | node1077 | node1079 | node1080 | node1083 | node1086 | node1087 | node1096 | node1115 | node1116 | node1222 | node1309 | node1328 | node1331 | node1342 | node1354 | node1386 | node1389 | node1393 | node1400 | node1413 | node1416 | node1428 | node1431 | node1436 | node1438 | node1445 | node1446 | node1448 | node1452 | node1453 | node1456 | node1459 | node1461 | node1475 | node1481 | node1490 | node1493 | node1497 | node1513 | node1521 | node1523 | node1524 | node1530 | node1540 | node1546 | node1552 | node1554 | node1562 | node1575 | node1587 | node1592 | node1597 | node1605 | node1607 | node1615 | node1622 | node1633 | node1637 | node1639 | node1640 | node1653 | node1673 | node1680 | node1776;
      result3 = node60 | node85 | node86 | node112 | node117 | node144 | node158 | node166 | node240 | node254 | node258 | node313 | node314 | node316 | node317 | node320 | node353 | node361 | node364 | node369 | node372 | node388 | node426 | node439 | node456 | node470 | node474 | node481 | node504 | node509 | node528 | node574 | node600 | node612 | node613 | node620 | node683 | node696 | node759 | node802 | node814 | node824 | node877 | node878 | node906 | node923 | node937 | node942 | node949 | node970 | node976 | node979 | node983 | node986 | node994 | node995 | node1017 | node1018 | node1026 | node1045 | node1052 | node1053 | node1055 | node1061 | node1076 | node1084 | node1094 | node1100 | node1104 | node1108 | node1109 | node1124 | node1125 | node1127 | node1131 | node1132 | node1134 | node1135 | node1139 | node1143 | node1146 | node1147 | node1150 | node1159 | node1198 | node1208 | node1221 | node1225 | node1245 | node1265 | node1268 | node1269 | node1275 | node1277 | node1285 | node1294 | node1301 | node1462 | node1551 | node1559 | node1600 | node1619 | node1631 | node1652 | node1669 | node1674 | node1679 | node1687 | node1690 | node1699 | node1715 | node1719 | node1726 | node1735 | node1738 | node1780 | node1785 | node1787 | node1803 | node1808;
      result4 = node10 | node11 | node14 | node18 | node32 | node36 | node58 | node82 | node125 | node126 | node131 | node136 | node140 | node161 | node164 | node174 | node178 | node189 | node191 | node284 | node291 | node349 | node356 | node362 | node381 | node397 | node443 | node465 | node542 | node555 | node577 | node598 | node604 | node648 | node669 | node692 | node695 | node700 | node702 | node708 | node710 | node714 | node715 | node718 | node727 | node730 | node734 | node738 | node744 | node745 | node766 | node813 | node820 | node823 | node829 | node853 | node862 | node863 | node868 | node901 | node1037 | node1290 | node1330 | node1335 | node1337 | node1358 | node1362 | node1385 | node1404 | node1432 | node1435 | node1496 | node1576 | node1583 | node1613 | node1661 | node1665 | node1686 | node1694 | node1718 | node1722 | node1732 | node1811;
      result5 = node33 | node44 | node57 | node71 | node98 | node101 | node104 | node109 | node116 | node152 | node154 | node160 | node167 | node177 | node185 | node229 | node249 | node287 | node292 | node294 | node299 | node300 | node302 | node321 | node329 | node331 | node347 | node350 | node403 | node410 | node415 | node480 | node487 | node493 | node502 | node505 | node518 | node567 | node569 | node573 | node581 | node582 | node584 | node585 | node622 | node632 | node660 | node674 | node681 | node723 | node724 | node726 | node737 | node741 | node751 | node754 | node771 | node780 | node787 | node788 | node803 | node816 | node817 | node859 | node874 | node891 | node905 | node926 | node930 | node934 | node952 | node955 | node984 | node987 | node991 | node998 | node999 | node1011 | node1014 | node1027 | node1111 | node1158 | node1165 | node1166 | node1168 | node1180 | node1183 | node1194 | node1201 | node1210 | node1228 | node1240 | node1246 | node1249 | node1255 | node1264 | node1271 | node1278 | node1293 | node1297 | node1298 | node1306 | node1312 | node1313 | node1348 | node1372 | node1465 | node1484 | node1544 | node1558 | node1677 | node1689 | node1706 | node1746 | node1760 | node1763 | node1781 | node1793 | node1800;
      result6 = node26 | node28 | node105 | node127 | node129 | node132 | node175 | node190 | node197 | node198 | node201 | node205 | node210 | node248 | node264 | node277 | node308 | node346 | node371 | node377 | node385 | node392 | node393 | node395 | node396 | node407 | node438 | node442 | node532 | node556 | node576 | node605 | node630 | node639 | node707 | node711 | node717 | node831 | node833 | node836 | node841 | node843 | node845 | node846 | node867 | node884 | node902 | node922 | node948 | node951 | node1177 | node1184 | node1190 | node1226 | node1238 | node1256 | node1281 | node1305 | node1316 | node1321 | node1324 | node1336 | node1347 | node1355 | node1357 | node1363 | node1382 | node1383 | node1392 | node1398 | node1421 | node1423 | node1424 | node1500 | node1508 | node1515 | node1528 | node1555 | node1569 | node1571 | node1572 | node1586 | node1590 | node1598 | node1608;
      result7 = node17 | node51 | node74 | node90 | node97 | node228 | node233 | node241 | node244 | node257 | node269 | node285 | node335 | node455 | node458 | node459 | node462 | node473 | node478 | node489 | node494 | node497 | node517 | node523 | node527 | node530 | node539 | node548 | node588 | node608 | node615 | node645 | node647 | node654 | node655 | node665 | node731 | node733 | node758 | node855 | node898 | node1604 | node1753 | node1770;
      result8 = node52 | node91 | node102 | node110 | node118 | node214 | node295 | node324 | node328 | node332 | node336 | node338 | node417 | node429 | node433 | node490 | node510 | node549 | node591 | node623 | node652 | node661 | node666 | node668 | node673 | node676 | node680 | node684 | node742 | node755 | node761 | node791 | node796 | node806 | node956 | node1001 | node1002 | node1010 | node1015 | node1046 | node1101 | node1103 | node1118 | node1119 | node1128 | node1140 | node1149 | node1161 | node1169 | node1176 | node1181 | node1195 | node1248 | node1272 | node1300 | node1315 | node1323 | node1341 | node1351 | node1373 | node1390 | node1397 | node1401 | node1405 | node1407 | node1408 | node1417 | node1420 | node1429 | node1439 | node1449 | node1455 | node1466 | node1468 | node1469 | node1474 | node1477 | node1478 | node1485 | node1492 | node1509 | node1512 | node1516 | node1531 | node1539 | node1543 | node1547 | node1561 | node1568 | node1578 | node1579 | node1584 | node1612 | node1616 | node1620 | node1623 | node1632 | node1636 | node1645 | node1648 | node1650 | node1658 | node1659 | node1662 | node1668 | node1676 | node1693 | node1695 | node1700 | node1702 | node1709 | node1710 | node1723 | node1725 | node1729 | node1731 | node1736 | node1739 | node1747 | node1749 | node1750 | node1754 | node1761 | node1764 | node1769 | node1772 | node1773 | node1777 | node1778 | node1788 | node1799 | node1802 | node1809 | node1816 | node1818 | node1819 | node1829 | node1830;
      result9 = node20 | node77 | node96 | node143 | node146 | node147 | node270 | node272 | node276 | node323 | node357 | node425 | node463 | node466 | node471 | node508 | node531 | node552 | node558 | node589 | node597 | node601 | node607 | node616 | node619 | node640 | node644 | node662 | node693 | node699 | node703 | node762 | node767 | node781 | node783 | node795 | node798 | node799 | node852 | node870 | node871 | node1056 | node1112 | node1235 | node1263 | node1291 | node1327 | node1414 | node1489 | node1703 | node1757 | node1792 | node1795 | node1812 | node1824;

      tree_5 = {result9, result8, result7, result6, result5, result4, result3, result2, result1, result0};
    end
  endfunction

  function [9:0] tree_6;
    input [783:0] pixel;

    reg node0_r;
    reg node0_l;
    reg node1_r;
    reg node1_l;
    reg node2_r;
    reg node2_l;
    reg node3_r;
    reg node3_l;
    reg node4_r;
    reg node4_l;
    reg node5_r;
    reg node5_l;
    reg node6_r;
    reg node6_l;
    reg node7_r;
    reg node7_l;
    reg node8_r;
    reg node8_l;
    reg node9_r;
    reg node9_l;
    reg node10;
    reg node11;
    reg node12_r;
    reg node12_l;
    reg node13;
    reg node14;
    reg node15_r;
    reg node15_l;
    reg node16_r;
    reg node16_l;
    reg node17;
    reg node18;
    reg node19_r;
    reg node19_l;
    reg node20;
    reg node21;
    reg node22_r;
    reg node22_l;
    reg node23_r;
    reg node23_l;
    reg node24_r;
    reg node24_l;
    reg node25;
    reg node26;
    reg node27_r;
    reg node27_l;
    reg node28;
    reg node29;
    reg node30_r;
    reg node30_l;
    reg node31_r;
    reg node31_l;
    reg node32;
    reg node33;
    reg node34_r;
    reg node34_l;
    reg node35;
    reg node36;
    reg node37_r;
    reg node37_l;
    reg node38_r;
    reg node38_l;
    reg node39_r;
    reg node39_l;
    reg node40_r;
    reg node40_l;
    reg node41;
    reg node42;
    reg node43_r;
    reg node43_l;
    reg node44;
    reg node45;
    reg node46_r;
    reg node46_l;
    reg node47_r;
    reg node47_l;
    reg node48;
    reg node49;
    reg node50_r;
    reg node50_l;
    reg node51;
    reg node52;
    reg node53_r;
    reg node53_l;
    reg node54_r;
    reg node54_l;
    reg node55_r;
    reg node55_l;
    reg node56;
    reg node57;
    reg node58_r;
    reg node58_l;
    reg node59;
    reg node60;
    reg node61_r;
    reg node61_l;
    reg node62_r;
    reg node62_l;
    reg node63;
    reg node64;
    reg node65_r;
    reg node65_l;
    reg node66;
    reg node67;
    reg node68_r;
    reg node68_l;
    reg node69_r;
    reg node69_l;
    reg node70_r;
    reg node70_l;
    reg node71_r;
    reg node71_l;
    reg node72_r;
    reg node72_l;
    reg node73;
    reg node74;
    reg node75_r;
    reg node75_l;
    reg node76;
    reg node77;
    reg node78_r;
    reg node78_l;
    reg node79_r;
    reg node79_l;
    reg node80;
    reg node81;
    reg node82_r;
    reg node82_l;
    reg node83;
    reg node84;
    reg node85_r;
    reg node85_l;
    reg node86_r;
    reg node86_l;
    reg node87_r;
    reg node87_l;
    reg node88;
    reg node89;
    reg node90_r;
    reg node90_l;
    reg node91;
    reg node92;
    reg node93_r;
    reg node93_l;
    reg node94_r;
    reg node94_l;
    reg node95;
    reg node96;
    reg node97_r;
    reg node97_l;
    reg node98;
    reg node99;
    reg node100_r;
    reg node100_l;
    reg node101_r;
    reg node101_l;
    reg node102_r;
    reg node102_l;
    reg node103_r;
    reg node103_l;
    reg node104;
    reg node105;
    reg node106_r;
    reg node106_l;
    reg node107;
    reg node108;
    reg node109_r;
    reg node109_l;
    reg node110_r;
    reg node110_l;
    reg node111;
    reg node112;
    reg node113_r;
    reg node113_l;
    reg node114;
    reg node115;
    reg node116_r;
    reg node116_l;
    reg node117_r;
    reg node117_l;
    reg node118_r;
    reg node118_l;
    reg node119;
    reg node120;
    reg node121_r;
    reg node121_l;
    reg node122;
    reg node123;
    reg node124_r;
    reg node124_l;
    reg node125_r;
    reg node125_l;
    reg node126;
    reg node127;
    reg node128_r;
    reg node128_l;
    reg node129;
    reg node130;
    reg node131_r;
    reg node131_l;
    reg node132_r;
    reg node132_l;
    reg node133_r;
    reg node133_l;
    reg node134_r;
    reg node134_l;
    reg node135_r;
    reg node135_l;
    reg node136_r;
    reg node136_l;
    reg node137;
    reg node138;
    reg node139_r;
    reg node139_l;
    reg node140;
    reg node141;
    reg node142_r;
    reg node142_l;
    reg node143_r;
    reg node143_l;
    reg node144;
    reg node145;
    reg node146_r;
    reg node146_l;
    reg node147;
    reg node148;
    reg node149_r;
    reg node149_l;
    reg node150_r;
    reg node150_l;
    reg node151_r;
    reg node151_l;
    reg node152;
    reg node153;
    reg node154_r;
    reg node154_l;
    reg node155;
    reg node156;
    reg node157_r;
    reg node157_l;
    reg node158_r;
    reg node158_l;
    reg node159;
    reg node160;
    reg node161_r;
    reg node161_l;
    reg node162;
    reg node163;
    reg node164_r;
    reg node164_l;
    reg node165_r;
    reg node165_l;
    reg node166_r;
    reg node166_l;
    reg node167_r;
    reg node167_l;
    reg node168;
    reg node169;
    reg node170;
    reg node171_r;
    reg node171_l;
    reg node172_r;
    reg node172_l;
    reg node173;
    reg node174;
    reg node175_r;
    reg node175_l;
    reg node176;
    reg node177;
    reg node178_r;
    reg node178_l;
    reg node179_r;
    reg node179_l;
    reg node180_r;
    reg node180_l;
    reg node181;
    reg node182;
    reg node183_r;
    reg node183_l;
    reg node184;
    reg node185;
    reg node186_r;
    reg node186_l;
    reg node187_r;
    reg node187_l;
    reg node188;
    reg node189;
    reg node190_r;
    reg node190_l;
    reg node191;
    reg node192;
    reg node193_r;
    reg node193_l;
    reg node194_r;
    reg node194_l;
    reg node195_r;
    reg node195_l;
    reg node196_r;
    reg node196_l;
    reg node197_r;
    reg node197_l;
    reg node198;
    reg node199;
    reg node200_r;
    reg node200_l;
    reg node201;
    reg node202;
    reg node203_r;
    reg node203_l;
    reg node204_r;
    reg node204_l;
    reg node205;
    reg node206;
    reg node207_r;
    reg node207_l;
    reg node208;
    reg node209;
    reg node210_r;
    reg node210_l;
    reg node211_r;
    reg node211_l;
    reg node212_r;
    reg node212_l;
    reg node213;
    reg node214;
    reg node215_r;
    reg node215_l;
    reg node216;
    reg node217;
    reg node218_r;
    reg node218_l;
    reg node219_r;
    reg node219_l;
    reg node220;
    reg node221;
    reg node222_r;
    reg node222_l;
    reg node223;
    reg node224;
    reg node225_r;
    reg node225_l;
    reg node226_r;
    reg node226_l;
    reg node227_r;
    reg node227_l;
    reg node228_r;
    reg node228_l;
    reg node229;
    reg node230;
    reg node231_r;
    reg node231_l;
    reg node232;
    reg node233;
    reg node234_r;
    reg node234_l;
    reg node235_r;
    reg node235_l;
    reg node236;
    reg node237;
    reg node238_r;
    reg node238_l;
    reg node239;
    reg node240;
    reg node241_r;
    reg node241_l;
    reg node242_r;
    reg node242_l;
    reg node243_r;
    reg node243_l;
    reg node244;
    reg node245;
    reg node246_r;
    reg node246_l;
    reg node247;
    reg node248;
    reg node249_r;
    reg node249_l;
    reg node250_r;
    reg node250_l;
    reg node251;
    reg node252;
    reg node253_r;
    reg node253_l;
    reg node254;
    reg node255;
    reg node256_r;
    reg node256_l;
    reg node257_r;
    reg node257_l;
    reg node258_r;
    reg node258_l;
    reg node259_r;
    reg node259_l;
    reg node260_r;
    reg node260_l;
    reg node261_r;
    reg node261_l;
    reg node262_r;
    reg node262_l;
    reg node263;
    reg node264;
    reg node265_r;
    reg node265_l;
    reg node266;
    reg node267;
    reg node268_r;
    reg node268_l;
    reg node269_r;
    reg node269_l;
    reg node270;
    reg node271;
    reg node272;
    reg node273_r;
    reg node273_l;
    reg node274_r;
    reg node274_l;
    reg node275_r;
    reg node275_l;
    reg node276;
    reg node277;
    reg node278_r;
    reg node278_l;
    reg node279;
    reg node280;
    reg node281_r;
    reg node281_l;
    reg node282_r;
    reg node282_l;
    reg node283;
    reg node284;
    reg node285_r;
    reg node285_l;
    reg node286;
    reg node287;
    reg node288_r;
    reg node288_l;
    reg node289_r;
    reg node289_l;
    reg node290_r;
    reg node290_l;
    reg node291_r;
    reg node291_l;
    reg node292;
    reg node293;
    reg node294_r;
    reg node294_l;
    reg node295;
    reg node296;
    reg node297_r;
    reg node297_l;
    reg node298_r;
    reg node298_l;
    reg node299;
    reg node300;
    reg node301_r;
    reg node301_l;
    reg node302;
    reg node303;
    reg node304_r;
    reg node304_l;
    reg node305_r;
    reg node305_l;
    reg node306_r;
    reg node306_l;
    reg node307;
    reg node308;
    reg node309;
    reg node310;
    reg node311_r;
    reg node311_l;
    reg node312_r;
    reg node312_l;
    reg node313_r;
    reg node313_l;
    reg node314_r;
    reg node314_l;
    reg node315_r;
    reg node315_l;
    reg node316;
    reg node317;
    reg node318_r;
    reg node318_l;
    reg node319;
    reg node320;
    reg node321_r;
    reg node321_l;
    reg node322_r;
    reg node322_l;
    reg node323;
    reg node324;
    reg node325_r;
    reg node325_l;
    reg node326;
    reg node327;
    reg node328_r;
    reg node328_l;
    reg node329_r;
    reg node329_l;
    reg node330;
    reg node331_r;
    reg node331_l;
    reg node332;
    reg node333;
    reg node334_r;
    reg node334_l;
    reg node335_r;
    reg node335_l;
    reg node336;
    reg node337;
    reg node338_r;
    reg node338_l;
    reg node339;
    reg node340;
    reg node341_r;
    reg node341_l;
    reg node342_r;
    reg node342_l;
    reg node343_r;
    reg node343_l;
    reg node344_r;
    reg node344_l;
    reg node345;
    reg node346;
    reg node347_r;
    reg node347_l;
    reg node348;
    reg node349;
    reg node350_r;
    reg node350_l;
    reg node351_r;
    reg node351_l;
    reg node352;
    reg node353;
    reg node354_r;
    reg node354_l;
    reg node355;
    reg node356;
    reg node357_r;
    reg node357_l;
    reg node358_r;
    reg node358_l;
    reg node359_r;
    reg node359_l;
    reg node360;
    reg node361;
    reg node362_r;
    reg node362_l;
    reg node363;
    reg node364;
    reg node365_r;
    reg node365_l;
    reg node366;
    reg node367_r;
    reg node367_l;
    reg node368;
    reg node369;
    reg node370_r;
    reg node370_l;
    reg node371_r;
    reg node371_l;
    reg node372_r;
    reg node372_l;
    reg node373_r;
    reg node373_l;
    reg node374_r;
    reg node374_l;
    reg node375_r;
    reg node375_l;
    reg node376;
    reg node377;
    reg node378_r;
    reg node378_l;
    reg node379;
    reg node380;
    reg node381_r;
    reg node381_l;
    reg node382_r;
    reg node382_l;
    reg node383;
    reg node384;
    reg node385_r;
    reg node385_l;
    reg node386;
    reg node387;
    reg node388_r;
    reg node388_l;
    reg node389_r;
    reg node389_l;
    reg node390_r;
    reg node390_l;
    reg node391;
    reg node392;
    reg node393_r;
    reg node393_l;
    reg node394;
    reg node395;
    reg node396_r;
    reg node396_l;
    reg node397_r;
    reg node397_l;
    reg node398;
    reg node399;
    reg node400_r;
    reg node400_l;
    reg node401;
    reg node402;
    reg node403_r;
    reg node403_l;
    reg node404_r;
    reg node404_l;
    reg node405_r;
    reg node405_l;
    reg node406_r;
    reg node406_l;
    reg node407;
    reg node408;
    reg node409_r;
    reg node409_l;
    reg node410;
    reg node411;
    reg node412_r;
    reg node412_l;
    reg node413_r;
    reg node413_l;
    reg node414;
    reg node415;
    reg node416_r;
    reg node416_l;
    reg node417;
    reg node418;
    reg node419_r;
    reg node419_l;
    reg node420_r;
    reg node420_l;
    reg node421_r;
    reg node421_l;
    reg node422;
    reg node423;
    reg node424_r;
    reg node424_l;
    reg node425;
    reg node426;
    reg node427_r;
    reg node427_l;
    reg node428_r;
    reg node428_l;
    reg node429;
    reg node430;
    reg node431_r;
    reg node431_l;
    reg node432;
    reg node433;
    reg node434_r;
    reg node434_l;
    reg node435_r;
    reg node435_l;
    reg node436_r;
    reg node436_l;
    reg node437_r;
    reg node437_l;
    reg node438_r;
    reg node438_l;
    reg node439;
    reg node440;
    reg node441_r;
    reg node441_l;
    reg node442;
    reg node443;
    reg node444_r;
    reg node444_l;
    reg node445_r;
    reg node445_l;
    reg node446;
    reg node447;
    reg node448_r;
    reg node448_l;
    reg node449;
    reg node450;
    reg node451_r;
    reg node451_l;
    reg node452_r;
    reg node452_l;
    reg node453_r;
    reg node453_l;
    reg node454;
    reg node455;
    reg node456_r;
    reg node456_l;
    reg node457;
    reg node458;
    reg node459_r;
    reg node459_l;
    reg node460_r;
    reg node460_l;
    reg node461;
    reg node462;
    reg node463;
    reg node464_r;
    reg node464_l;
    reg node465_r;
    reg node465_l;
    reg node466_r;
    reg node466_l;
    reg node467_r;
    reg node467_l;
    reg node468;
    reg node469;
    reg node470_r;
    reg node470_l;
    reg node471;
    reg node472;
    reg node473_r;
    reg node473_l;
    reg node474_r;
    reg node474_l;
    reg node475;
    reg node476;
    reg node477_r;
    reg node477_l;
    reg node478;
    reg node479;
    reg node480_r;
    reg node480_l;
    reg node481_r;
    reg node481_l;
    reg node482_r;
    reg node482_l;
    reg node483;
    reg node484;
    reg node485;
    reg node486_r;
    reg node486_l;
    reg node487_r;
    reg node487_l;
    reg node488;
    reg node489;
    reg node490_r;
    reg node490_l;
    reg node491;
    reg node492;
    reg node493_r;
    reg node493_l;
    reg node494_r;
    reg node494_l;
    reg node495_r;
    reg node495_l;
    reg node496_r;
    reg node496_l;
    reg node497_r;
    reg node497_l;
    reg node498_r;
    reg node498_l;
    reg node499_r;
    reg node499_l;
    reg node500_r;
    reg node500_l;
    reg node501;
    reg node502;
    reg node503_r;
    reg node503_l;
    reg node504;
    reg node505;
    reg node506_r;
    reg node506_l;
    reg node507_r;
    reg node507_l;
    reg node508;
    reg node509;
    reg node510;
    reg node511_r;
    reg node511_l;
    reg node512_r;
    reg node512_l;
    reg node513_r;
    reg node513_l;
    reg node514;
    reg node515;
    reg node516_r;
    reg node516_l;
    reg node517;
    reg node518;
    reg node519_r;
    reg node519_l;
    reg node520_r;
    reg node520_l;
    reg node521;
    reg node522;
    reg node523_r;
    reg node523_l;
    reg node524;
    reg node525;
    reg node526_r;
    reg node526_l;
    reg node527_r;
    reg node527_l;
    reg node528_r;
    reg node528_l;
    reg node529_r;
    reg node529_l;
    reg node530;
    reg node531;
    reg node532_r;
    reg node532_l;
    reg node533;
    reg node534;
    reg node535_r;
    reg node535_l;
    reg node536;
    reg node537;
    reg node538_r;
    reg node538_l;
    reg node539_r;
    reg node539_l;
    reg node540;
    reg node541_r;
    reg node541_l;
    reg node542;
    reg node543;
    reg node544;
    reg node545_r;
    reg node545_l;
    reg node546_r;
    reg node546_l;
    reg node547_r;
    reg node547_l;
    reg node548_r;
    reg node548_l;
    reg node549_r;
    reg node549_l;
    reg node550;
    reg node551;
    reg node552_r;
    reg node552_l;
    reg node553;
    reg node554;
    reg node555_r;
    reg node555_l;
    reg node556;
    reg node557_r;
    reg node557_l;
    reg node558;
    reg node559;
    reg node560_r;
    reg node560_l;
    reg node561_r;
    reg node561_l;
    reg node562_r;
    reg node562_l;
    reg node563;
    reg node564;
    reg node565_r;
    reg node565_l;
    reg node566;
    reg node567;
    reg node568_r;
    reg node568_l;
    reg node569_r;
    reg node569_l;
    reg node570;
    reg node571;
    reg node572;
    reg node573_r;
    reg node573_l;
    reg node574_r;
    reg node574_l;
    reg node575_r;
    reg node575_l;
    reg node576_r;
    reg node576_l;
    reg node577;
    reg node578;
    reg node579_r;
    reg node579_l;
    reg node580;
    reg node581;
    reg node582_r;
    reg node582_l;
    reg node583_r;
    reg node583_l;
    reg node584;
    reg node585;
    reg node586_r;
    reg node586_l;
    reg node587;
    reg node588;
    reg node589_r;
    reg node589_l;
    reg node590_r;
    reg node590_l;
    reg node591_r;
    reg node591_l;
    reg node592;
    reg node593;
    reg node594_r;
    reg node594_l;
    reg node595;
    reg node596;
    reg node597_r;
    reg node597_l;
    reg node598_r;
    reg node598_l;
    reg node599;
    reg node600;
    reg node601_r;
    reg node601_l;
    reg node602;
    reg node603;
    reg node604_r;
    reg node604_l;
    reg node605_r;
    reg node605_l;
    reg node606_r;
    reg node606_l;
    reg node607_r;
    reg node607_l;
    reg node608_r;
    reg node608_l;
    reg node609_r;
    reg node609_l;
    reg node610;
    reg node611;
    reg node612;
    reg node613_r;
    reg node613_l;
    reg node614_r;
    reg node614_l;
    reg node615;
    reg node616;
    reg node617_r;
    reg node617_l;
    reg node618;
    reg node619;
    reg node620_r;
    reg node620_l;
    reg node621_r;
    reg node621_l;
    reg node622;
    reg node623_r;
    reg node623_l;
    reg node624;
    reg node625;
    reg node626_r;
    reg node626_l;
    reg node627;
    reg node628;
    reg node629_r;
    reg node629_l;
    reg node630_r;
    reg node630_l;
    reg node631_r;
    reg node631_l;
    reg node632_r;
    reg node632_l;
    reg node633;
    reg node634;
    reg node635_r;
    reg node635_l;
    reg node636;
    reg node637;
    reg node638_r;
    reg node638_l;
    reg node639_r;
    reg node639_l;
    reg node640;
    reg node641;
    reg node642_r;
    reg node642_l;
    reg node643;
    reg node644;
    reg node645_r;
    reg node645_l;
    reg node646;
    reg node647_r;
    reg node647_l;
    reg node648;
    reg node649;
    reg node650_r;
    reg node650_l;
    reg node651;
    reg node652_r;
    reg node652_l;
    reg node653_r;
    reg node653_l;
    reg node654;
    reg node655_r;
    reg node655_l;
    reg node656;
    reg node657;
    reg node658_r;
    reg node658_l;
    reg node659;
    reg node660_r;
    reg node660_l;
    reg node661;
    reg node662;
    reg node663_r;
    reg node663_l;
    reg node664_r;
    reg node664_l;
    reg node665_r;
    reg node665_l;
    reg node666_r;
    reg node666_l;
    reg node667_r;
    reg node667_l;
    reg node668_r;
    reg node668_l;
    reg node669_r;
    reg node669_l;
    reg node670;
    reg node671;
    reg node672_r;
    reg node672_l;
    reg node673;
    reg node674;
    reg node675;
    reg node676;
    reg node677_r;
    reg node677_l;
    reg node678_r;
    reg node678_l;
    reg node679_r;
    reg node679_l;
    reg node680_r;
    reg node680_l;
    reg node681;
    reg node682;
    reg node683;
    reg node684;
    reg node685_r;
    reg node685_l;
    reg node686;
    reg node687;
    reg node688_r;
    reg node688_l;
    reg node689_r;
    reg node689_l;
    reg node690_r;
    reg node690_l;
    reg node691_r;
    reg node691_l;
    reg node692_r;
    reg node692_l;
    reg node693;
    reg node694;
    reg node695_r;
    reg node695_l;
    reg node696;
    reg node697;
    reg node698_r;
    reg node698_l;
    reg node699;
    reg node700_r;
    reg node700_l;
    reg node701;
    reg node702;
    reg node703_r;
    reg node703_l;
    reg node704_r;
    reg node704_l;
    reg node705;
    reg node706;
    reg node707_r;
    reg node707_l;
    reg node708;
    reg node709;
    reg node710_r;
    reg node710_l;
    reg node711_r;
    reg node711_l;
    reg node712_r;
    reg node712_l;
    reg node713_r;
    reg node713_l;
    reg node714;
    reg node715;
    reg node716;
    reg node717_r;
    reg node717_l;
    reg node718;
    reg node719_r;
    reg node719_l;
    reg node720;
    reg node721;
    reg node722_r;
    reg node722_l;
    reg node723_r;
    reg node723_l;
    reg node724;
    reg node725;
    reg node726_r;
    reg node726_l;
    reg node727_r;
    reg node727_l;
    reg node728;
    reg node729;
    reg node730;
    reg node731_r;
    reg node731_l;
    reg node732_r;
    reg node732_l;
    reg node733_r;
    reg node733_l;
    reg node734_r;
    reg node734_l;
    reg node735_r;
    reg node735_l;
    reg node736_r;
    reg node736_l;
    reg node737;
    reg node738;
    reg node739_r;
    reg node739_l;
    reg node740;
    reg node741;
    reg node742_r;
    reg node742_l;
    reg node743_r;
    reg node743_l;
    reg node744;
    reg node745;
    reg node746_r;
    reg node746_l;
    reg node747;
    reg node748;
    reg node749_r;
    reg node749_l;
    reg node750_r;
    reg node750_l;
    reg node751_r;
    reg node751_l;
    reg node752;
    reg node753;
    reg node754_r;
    reg node754_l;
    reg node755;
    reg node756;
    reg node757_r;
    reg node757_l;
    reg node758_r;
    reg node758_l;
    reg node759;
    reg node760;
    reg node761_r;
    reg node761_l;
    reg node762;
    reg node763;
    reg node764_r;
    reg node764_l;
    reg node765_r;
    reg node765_l;
    reg node766_r;
    reg node766_l;
    reg node767_r;
    reg node767_l;
    reg node768;
    reg node769;
    reg node770;
    reg node771;
    reg node772;
    reg node773_r;
    reg node773_l;
    reg node774_r;
    reg node774_l;
    reg node775_r;
    reg node775_l;
    reg node776_r;
    reg node776_l;
    reg node777_r;
    reg node777_l;
    reg node778;
    reg node779;
    reg node780;
    reg node781_r;
    reg node781_l;
    reg node782_r;
    reg node782_l;
    reg node783;
    reg node784;
    reg node785_r;
    reg node785_l;
    reg node786;
    reg node787;
    reg node788_r;
    reg node788_l;
    reg node789_r;
    reg node789_l;
    reg node790_r;
    reg node790_l;
    reg node791;
    reg node792;
    reg node793_r;
    reg node793_l;
    reg node794;
    reg node795;
    reg node796_r;
    reg node796_l;
    reg node797_r;
    reg node797_l;
    reg node798;
    reg node799;
    reg node800_r;
    reg node800_l;
    reg node801;
    reg node802;
    reg node803_r;
    reg node803_l;
    reg node804_r;
    reg node804_l;
    reg node805_r;
    reg node805_l;
    reg node806_r;
    reg node806_l;
    reg node807;
    reg node808;
    reg node809_r;
    reg node809_l;
    reg node810;
    reg node811;
    reg node812_r;
    reg node812_l;
    reg node813_r;
    reg node813_l;
    reg node814;
    reg node815;
    reg node816_r;
    reg node816_l;
    reg node817;
    reg node818;
    reg node819_r;
    reg node819_l;
    reg node820_r;
    reg node820_l;
    reg node821_r;
    reg node821_l;
    reg node822;
    reg node823;
    reg node824_r;
    reg node824_l;
    reg node825;
    reg node826;
    reg node827_r;
    reg node827_l;
    reg node828_r;
    reg node828_l;
    reg node829;
    reg node830;
    reg node831_r;
    reg node831_l;
    reg node832;
    reg node833;
    reg node834_r;
    reg node834_l;
    reg node835_r;
    reg node835_l;
    reg node836_r;
    reg node836_l;
    reg node837_r;
    reg node837_l;
    reg node838_r;
    reg node838_l;
    reg node839_r;
    reg node839_l;
    reg node840_r;
    reg node840_l;
    reg node841_r;
    reg node841_l;
    reg node842_r;
    reg node842_l;
    reg node843;
    reg node844;
    reg node845_r;
    reg node845_l;
    reg node846;
    reg node847;
    reg node848_r;
    reg node848_l;
    reg node849_r;
    reg node849_l;
    reg node850;
    reg node851;
    reg node852_r;
    reg node852_l;
    reg node853;
    reg node854;
    reg node855_r;
    reg node855_l;
    reg node856_r;
    reg node856_l;
    reg node857_r;
    reg node857_l;
    reg node858;
    reg node859;
    reg node860_r;
    reg node860_l;
    reg node861;
    reg node862;
    reg node863_r;
    reg node863_l;
    reg node864_r;
    reg node864_l;
    reg node865;
    reg node866;
    reg node867_r;
    reg node867_l;
    reg node868;
    reg node869;
    reg node870_r;
    reg node870_l;
    reg node871_r;
    reg node871_l;
    reg node872_r;
    reg node872_l;
    reg node873_r;
    reg node873_l;
    reg node874;
    reg node875;
    reg node876_r;
    reg node876_l;
    reg node877;
    reg node878;
    reg node879_r;
    reg node879_l;
    reg node880_r;
    reg node880_l;
    reg node881;
    reg node882;
    reg node883_r;
    reg node883_l;
    reg node884;
    reg node885;
    reg node886_r;
    reg node886_l;
    reg node887_r;
    reg node887_l;
    reg node888;
    reg node889;
    reg node890_r;
    reg node890_l;
    reg node891_r;
    reg node891_l;
    reg node892;
    reg node893;
    reg node894;
    reg node895_r;
    reg node895_l;
    reg node896_r;
    reg node896_l;
    reg node897_r;
    reg node897_l;
    reg node898_r;
    reg node898_l;
    reg node899_r;
    reg node899_l;
    reg node900;
    reg node901;
    reg node902_r;
    reg node902_l;
    reg node903;
    reg node904;
    reg node905_r;
    reg node905_l;
    reg node906_r;
    reg node906_l;
    reg node907;
    reg node908;
    reg node909_r;
    reg node909_l;
    reg node910;
    reg node911;
    reg node912_r;
    reg node912_l;
    reg node913_r;
    reg node913_l;
    reg node914_r;
    reg node914_l;
    reg node915;
    reg node916;
    reg node917_r;
    reg node917_l;
    reg node918;
    reg node919;
    reg node920_r;
    reg node920_l;
    reg node921_r;
    reg node921_l;
    reg node922;
    reg node923;
    reg node924;
    reg node925_r;
    reg node925_l;
    reg node926_r;
    reg node926_l;
    reg node927_r;
    reg node927_l;
    reg node928_r;
    reg node928_l;
    reg node929;
    reg node930;
    reg node931_r;
    reg node931_l;
    reg node932;
    reg node933;
    reg node934_r;
    reg node934_l;
    reg node935_r;
    reg node935_l;
    reg node936;
    reg node937;
    reg node938;
    reg node939_r;
    reg node939_l;
    reg node940_r;
    reg node940_l;
    reg node941_r;
    reg node941_l;
    reg node942;
    reg node943;
    reg node944_r;
    reg node944_l;
    reg node945;
    reg node946;
    reg node947_r;
    reg node947_l;
    reg node948;
    reg node949_r;
    reg node949_l;
    reg node950;
    reg node951;
    reg node952_r;
    reg node952_l;
    reg node953_r;
    reg node953_l;
    reg node954_r;
    reg node954_l;
    reg node955_r;
    reg node955_l;
    reg node956_r;
    reg node956_l;
    reg node957_r;
    reg node957_l;
    reg node958;
    reg node959;
    reg node960_r;
    reg node960_l;
    reg node961;
    reg node962;
    reg node963_r;
    reg node963_l;
    reg node964;
    reg node965_r;
    reg node965_l;
    reg node966;
    reg node967;
    reg node968_r;
    reg node968_l;
    reg node969_r;
    reg node969_l;
    reg node970_r;
    reg node970_l;
    reg node971;
    reg node972;
    reg node973_r;
    reg node973_l;
    reg node974;
    reg node975;
    reg node976_r;
    reg node976_l;
    reg node977_r;
    reg node977_l;
    reg node978;
    reg node979;
    reg node980_r;
    reg node980_l;
    reg node981;
    reg node982;
    reg node983_r;
    reg node983_l;
    reg node984_r;
    reg node984_l;
    reg node985_r;
    reg node985_l;
    reg node986_r;
    reg node986_l;
    reg node987;
    reg node988;
    reg node989_r;
    reg node989_l;
    reg node990;
    reg node991;
    reg node992_r;
    reg node992_l;
    reg node993_r;
    reg node993_l;
    reg node994;
    reg node995;
    reg node996_r;
    reg node996_l;
    reg node997;
    reg node998;
    reg node999_r;
    reg node999_l;
    reg node1000_r;
    reg node1000_l;
    reg node1001_r;
    reg node1001_l;
    reg node1002;
    reg node1003;
    reg node1004_r;
    reg node1004_l;
    reg node1005;
    reg node1006;
    reg node1007_r;
    reg node1007_l;
    reg node1008_r;
    reg node1008_l;
    reg node1009;
    reg node1010;
    reg node1011_r;
    reg node1011_l;
    reg node1012;
    reg node1013;
    reg node1014_r;
    reg node1014_l;
    reg node1015_r;
    reg node1015_l;
    reg node1016_r;
    reg node1016_l;
    reg node1017_r;
    reg node1017_l;
    reg node1018_r;
    reg node1018_l;
    reg node1019;
    reg node1020;
    reg node1021_r;
    reg node1021_l;
    reg node1022;
    reg node1023;
    reg node1024_r;
    reg node1024_l;
    reg node1025_r;
    reg node1025_l;
    reg node1026;
    reg node1027;
    reg node1028_r;
    reg node1028_l;
    reg node1029;
    reg node1030;
    reg node1031_r;
    reg node1031_l;
    reg node1032_r;
    reg node1032_l;
    reg node1033_r;
    reg node1033_l;
    reg node1034;
    reg node1035;
    reg node1036_r;
    reg node1036_l;
    reg node1037;
    reg node1038;
    reg node1039_r;
    reg node1039_l;
    reg node1040_r;
    reg node1040_l;
    reg node1041;
    reg node1042;
    reg node1043_r;
    reg node1043_l;
    reg node1044;
    reg node1045;
    reg node1046_r;
    reg node1046_l;
    reg node1047_r;
    reg node1047_l;
    reg node1048_r;
    reg node1048_l;
    reg node1049_r;
    reg node1049_l;
    reg node1050;
    reg node1051;
    reg node1052_r;
    reg node1052_l;
    reg node1053;
    reg node1054;
    reg node1055_r;
    reg node1055_l;
    reg node1056_r;
    reg node1056_l;
    reg node1057;
    reg node1058;
    reg node1059_r;
    reg node1059_l;
    reg node1060;
    reg node1061;
    reg node1062_r;
    reg node1062_l;
    reg node1063_r;
    reg node1063_l;
    reg node1064_r;
    reg node1064_l;
    reg node1065;
    reg node1066;
    reg node1067_r;
    reg node1067_l;
    reg node1068;
    reg node1069;
    reg node1070_r;
    reg node1070_l;
    reg node1071_r;
    reg node1071_l;
    reg node1072;
    reg node1073;
    reg node1074_r;
    reg node1074_l;
    reg node1075;
    reg node1076;
    reg node1077_r;
    reg node1077_l;
    reg node1078_r;
    reg node1078_l;
    reg node1079_r;
    reg node1079_l;
    reg node1080_r;
    reg node1080_l;
    reg node1081_r;
    reg node1081_l;
    reg node1082_r;
    reg node1082_l;
    reg node1083_r;
    reg node1083_l;
    reg node1084;
    reg node1085;
    reg node1086_r;
    reg node1086_l;
    reg node1087;
    reg node1088;
    reg node1089_r;
    reg node1089_l;
    reg node1090_r;
    reg node1090_l;
    reg node1091;
    reg node1092;
    reg node1093_r;
    reg node1093_l;
    reg node1094;
    reg node1095;
    reg node1096_r;
    reg node1096_l;
    reg node1097_r;
    reg node1097_l;
    reg node1098_r;
    reg node1098_l;
    reg node1099;
    reg node1100;
    reg node1101_r;
    reg node1101_l;
    reg node1102;
    reg node1103;
    reg node1104_r;
    reg node1104_l;
    reg node1105_r;
    reg node1105_l;
    reg node1106;
    reg node1107;
    reg node1108;
    reg node1109_r;
    reg node1109_l;
    reg node1110_r;
    reg node1110_l;
    reg node1111_r;
    reg node1111_l;
    reg node1112_r;
    reg node1112_l;
    reg node1113;
    reg node1114;
    reg node1115_r;
    reg node1115_l;
    reg node1116;
    reg node1117;
    reg node1118_r;
    reg node1118_l;
    reg node1119_r;
    reg node1119_l;
    reg node1120;
    reg node1121;
    reg node1122_r;
    reg node1122_l;
    reg node1123;
    reg node1124;
    reg node1125_r;
    reg node1125_l;
    reg node1126_r;
    reg node1126_l;
    reg node1127_r;
    reg node1127_l;
    reg node1128;
    reg node1129;
    reg node1130_r;
    reg node1130_l;
    reg node1131;
    reg node1132;
    reg node1133_r;
    reg node1133_l;
    reg node1134_r;
    reg node1134_l;
    reg node1135;
    reg node1136;
    reg node1137;
    reg node1138_r;
    reg node1138_l;
    reg node1139_r;
    reg node1139_l;
    reg node1140_r;
    reg node1140_l;
    reg node1141_r;
    reg node1141_l;
    reg node1142_r;
    reg node1142_l;
    reg node1143;
    reg node1144;
    reg node1145_r;
    reg node1145_l;
    reg node1146;
    reg node1147;
    reg node1148;
    reg node1149_r;
    reg node1149_l;
    reg node1150_r;
    reg node1150_l;
    reg node1151;
    reg node1152;
    reg node1153_r;
    reg node1153_l;
    reg node1154_r;
    reg node1154_l;
    reg node1155;
    reg node1156;
    reg node1157_r;
    reg node1157_l;
    reg node1158;
    reg node1159;
    reg node1160_r;
    reg node1160_l;
    reg node1161_r;
    reg node1161_l;
    reg node1162_r;
    reg node1162_l;
    reg node1163_r;
    reg node1163_l;
    reg node1164;
    reg node1165;
    reg node1166_r;
    reg node1166_l;
    reg node1167;
    reg node1168;
    reg node1169_r;
    reg node1169_l;
    reg node1170_r;
    reg node1170_l;
    reg node1171;
    reg node1172;
    reg node1173_r;
    reg node1173_l;
    reg node1174;
    reg node1175;
    reg node1176_r;
    reg node1176_l;
    reg node1177_r;
    reg node1177_l;
    reg node1178_r;
    reg node1178_l;
    reg node1179;
    reg node1180;
    reg node1181;
    reg node1182_r;
    reg node1182_l;
    reg node1183_r;
    reg node1183_l;
    reg node1184;
    reg node1185;
    reg node1186_r;
    reg node1186_l;
    reg node1187;
    reg node1188;
    reg node1189_r;
    reg node1189_l;
    reg node1190_r;
    reg node1190_l;
    reg node1191_r;
    reg node1191_l;
    reg node1192_r;
    reg node1192_l;
    reg node1193_r;
    reg node1193_l;
    reg node1194_r;
    reg node1194_l;
    reg node1195;
    reg node1196;
    reg node1197_r;
    reg node1197_l;
    reg node1198;
    reg node1199;
    reg node1200_r;
    reg node1200_l;
    reg node1201_r;
    reg node1201_l;
    reg node1202;
    reg node1203;
    reg node1204_r;
    reg node1204_l;
    reg node1205;
    reg node1206;
    reg node1207_r;
    reg node1207_l;
    reg node1208_r;
    reg node1208_l;
    reg node1209_r;
    reg node1209_l;
    reg node1210;
    reg node1211;
    reg node1212_r;
    reg node1212_l;
    reg node1213;
    reg node1214;
    reg node1215_r;
    reg node1215_l;
    reg node1216_r;
    reg node1216_l;
    reg node1217;
    reg node1218;
    reg node1219_r;
    reg node1219_l;
    reg node1220;
    reg node1221;
    reg node1222_r;
    reg node1222_l;
    reg node1223_r;
    reg node1223_l;
    reg node1224_r;
    reg node1224_l;
    reg node1225_r;
    reg node1225_l;
    reg node1226;
    reg node1227;
    reg node1228_r;
    reg node1228_l;
    reg node1229;
    reg node1230;
    reg node1231_r;
    reg node1231_l;
    reg node1232;
    reg node1233;
    reg node1234_r;
    reg node1234_l;
    reg node1235_r;
    reg node1235_l;
    reg node1236;
    reg node1237_r;
    reg node1237_l;
    reg node1238;
    reg node1239;
    reg node1240;
    reg node1241_r;
    reg node1241_l;
    reg node1242_r;
    reg node1242_l;
    reg node1243_r;
    reg node1243_l;
    reg node1244_r;
    reg node1244_l;
    reg node1245_r;
    reg node1245_l;
    reg node1246;
    reg node1247;
    reg node1248_r;
    reg node1248_l;
    reg node1249;
    reg node1250;
    reg node1251_r;
    reg node1251_l;
    reg node1252_r;
    reg node1252_l;
    reg node1253;
    reg node1254;
    reg node1255_r;
    reg node1255_l;
    reg node1256;
    reg node1257;
    reg node1258_r;
    reg node1258_l;
    reg node1259_r;
    reg node1259_l;
    reg node1260_r;
    reg node1260_l;
    reg node1261;
    reg node1262;
    reg node1263;
    reg node1264_r;
    reg node1264_l;
    reg node1265_r;
    reg node1265_l;
    reg node1266;
    reg node1267;
    reg node1268_r;
    reg node1268_l;
    reg node1269;
    reg node1270;
    reg node1271_r;
    reg node1271_l;
    reg node1272_r;
    reg node1272_l;
    reg node1273;
    reg node1274;
    reg node1275_r;
    reg node1275_l;
    reg node1276_r;
    reg node1276_l;
    reg node1277;
    reg node1278_r;
    reg node1278_l;
    reg node1279;
    reg node1280;
    reg node1281_r;
    reg node1281_l;
    reg node1282_r;
    reg node1282_l;
    reg node1283;
    reg node1284;
    reg node1285_r;
    reg node1285_l;
    reg node1286;
    reg node1287;
    reg node1288_r;
    reg node1288_l;
    reg node1289_r;
    reg node1289_l;
    reg node1290_r;
    reg node1290_l;
    reg node1291_r;
    reg node1291_l;
    reg node1292_r;
    reg node1292_l;
    reg node1293_r;
    reg node1293_l;
    reg node1294_r;
    reg node1294_l;
    reg node1295_r;
    reg node1295_l;
    reg node1296;
    reg node1297;
    reg node1298;
    reg node1299_r;
    reg node1299_l;
    reg node1300_r;
    reg node1300_l;
    reg node1301;
    reg node1302;
    reg node1303_r;
    reg node1303_l;
    reg node1304;
    reg node1305;
    reg node1306_r;
    reg node1306_l;
    reg node1307_r;
    reg node1307_l;
    reg node1308_r;
    reg node1308_l;
    reg node1309;
    reg node1310;
    reg node1311_r;
    reg node1311_l;
    reg node1312;
    reg node1313;
    reg node1314_r;
    reg node1314_l;
    reg node1315_r;
    reg node1315_l;
    reg node1316;
    reg node1317;
    reg node1318_r;
    reg node1318_l;
    reg node1319;
    reg node1320;
    reg node1321_r;
    reg node1321_l;
    reg node1322_r;
    reg node1322_l;
    reg node1323_r;
    reg node1323_l;
    reg node1324_r;
    reg node1324_l;
    reg node1325;
    reg node1326;
    reg node1327_r;
    reg node1327_l;
    reg node1328;
    reg node1329;
    reg node1330_r;
    reg node1330_l;
    reg node1331_r;
    reg node1331_l;
    reg node1332;
    reg node1333;
    reg node1334_r;
    reg node1334_l;
    reg node1335;
    reg node1336;
    reg node1337_r;
    reg node1337_l;
    reg node1338_r;
    reg node1338_l;
    reg node1339_r;
    reg node1339_l;
    reg node1340;
    reg node1341;
    reg node1342_r;
    reg node1342_l;
    reg node1343;
    reg node1344;
    reg node1345_r;
    reg node1345_l;
    reg node1346_r;
    reg node1346_l;
    reg node1347;
    reg node1348;
    reg node1349_r;
    reg node1349_l;
    reg node1350;
    reg node1351;
    reg node1352_r;
    reg node1352_l;
    reg node1353_r;
    reg node1353_l;
    reg node1354_r;
    reg node1354_l;
    reg node1355_r;
    reg node1355_l;
    reg node1356_r;
    reg node1356_l;
    reg node1357;
    reg node1358;
    reg node1359_r;
    reg node1359_l;
    reg node1360;
    reg node1361;
    reg node1362_r;
    reg node1362_l;
    reg node1363_r;
    reg node1363_l;
    reg node1364;
    reg node1365;
    reg node1366_r;
    reg node1366_l;
    reg node1367;
    reg node1368;
    reg node1369_r;
    reg node1369_l;
    reg node1370_r;
    reg node1370_l;
    reg node1371_r;
    reg node1371_l;
    reg node1372;
    reg node1373;
    reg node1374_r;
    reg node1374_l;
    reg node1375;
    reg node1376;
    reg node1377_r;
    reg node1377_l;
    reg node1378_r;
    reg node1378_l;
    reg node1379;
    reg node1380;
    reg node1381_r;
    reg node1381_l;
    reg node1382;
    reg node1383;
    reg node1384_r;
    reg node1384_l;
    reg node1385_r;
    reg node1385_l;
    reg node1386_r;
    reg node1386_l;
    reg node1387_r;
    reg node1387_l;
    reg node1388;
    reg node1389;
    reg node1390_r;
    reg node1390_l;
    reg node1391;
    reg node1392;
    reg node1393_r;
    reg node1393_l;
    reg node1394;
    reg node1395_r;
    reg node1395_l;
    reg node1396;
    reg node1397;
    reg node1398_r;
    reg node1398_l;
    reg node1399_r;
    reg node1399_l;
    reg node1400_r;
    reg node1400_l;
    reg node1401;
    reg node1402;
    reg node1403_r;
    reg node1403_l;
    reg node1404;
    reg node1405;
    reg node1406_r;
    reg node1406_l;
    reg node1407_r;
    reg node1407_l;
    reg node1408;
    reg node1409;
    reg node1410_r;
    reg node1410_l;
    reg node1411;
    reg node1412;
    reg node1413_r;
    reg node1413_l;
    reg node1414_r;
    reg node1414_l;
    reg node1415_r;
    reg node1415_l;
    reg node1416_r;
    reg node1416_l;
    reg node1417_r;
    reg node1417_l;
    reg node1418_r;
    reg node1418_l;
    reg node1419;
    reg node1420;
    reg node1421_r;
    reg node1421_l;
    reg node1422;
    reg node1423;
    reg node1424_r;
    reg node1424_l;
    reg node1425_r;
    reg node1425_l;
    reg node1426;
    reg node1427;
    reg node1428;
    reg node1429_r;
    reg node1429_l;
    reg node1430_r;
    reg node1430_l;
    reg node1431;
    reg node1432;
    reg node1433_r;
    reg node1433_l;
    reg node1434;
    reg node1435_r;
    reg node1435_l;
    reg node1436;
    reg node1437;
    reg node1438_r;
    reg node1438_l;
    reg node1439;
    reg node1440;
    reg node1441_r;
    reg node1441_l;
    reg node1442_r;
    reg node1442_l;
    reg node1443_r;
    reg node1443_l;
    reg node1444_r;
    reg node1444_l;
    reg node1445_r;
    reg node1445_l;
    reg node1446;
    reg node1447;
    reg node1448;
    reg node1449_r;
    reg node1449_l;
    reg node1450_r;
    reg node1450_l;
    reg node1451;
    reg node1452;
    reg node1453;
    reg node1454_r;
    reg node1454_l;
    reg node1455_r;
    reg node1455_l;
    reg node1456;
    reg node1457;
    reg node1458;
    reg node1459_r;
    reg node1459_l;
    reg node1460_r;
    reg node1460_l;
    reg node1461_r;
    reg node1461_l;
    reg node1462;
    reg node1463;
    reg node1464;
    reg node1465_r;
    reg node1465_l;
    reg node1466;
    reg node1467_r;
    reg node1467_l;
    reg node1468;
    reg node1469;
    reg node1470_r;
    reg node1470_l;
    reg node1471_r;
    reg node1471_l;
    reg node1472_r;
    reg node1472_l;
    reg node1473_r;
    reg node1473_l;
    reg node1474_r;
    reg node1474_l;
    reg node1475_r;
    reg node1475_l;
    reg node1476_r;
    reg node1476_l;
    reg node1477;
    reg node1478;
    reg node1479_r;
    reg node1479_l;
    reg node1480;
    reg node1481;
    reg node1482_r;
    reg node1482_l;
    reg node1483_r;
    reg node1483_l;
    reg node1484;
    reg node1485;
    reg node1486_r;
    reg node1486_l;
    reg node1487;
    reg node1488;
    reg node1489_r;
    reg node1489_l;
    reg node1490_r;
    reg node1490_l;
    reg node1491_r;
    reg node1491_l;
    reg node1492;
    reg node1493;
    reg node1494_r;
    reg node1494_l;
    reg node1495;
    reg node1496;
    reg node1497_r;
    reg node1497_l;
    reg node1498_r;
    reg node1498_l;
    reg node1499;
    reg node1500;
    reg node1501_r;
    reg node1501_l;
    reg node1502;
    reg node1503;
    reg node1504_r;
    reg node1504_l;
    reg node1505_r;
    reg node1505_l;
    reg node1506_r;
    reg node1506_l;
    reg node1507_r;
    reg node1507_l;
    reg node1508;
    reg node1509;
    reg node1510_r;
    reg node1510_l;
    reg node1511;
    reg node1512;
    reg node1513_r;
    reg node1513_l;
    reg node1514_r;
    reg node1514_l;
    reg node1515;
    reg node1516;
    reg node1517_r;
    reg node1517_l;
    reg node1518;
    reg node1519;
    reg node1520_r;
    reg node1520_l;
    reg node1521_r;
    reg node1521_l;
    reg node1522_r;
    reg node1522_l;
    reg node1523;
    reg node1524;
    reg node1525_r;
    reg node1525_l;
    reg node1526;
    reg node1527;
    reg node1528_r;
    reg node1528_l;
    reg node1529_r;
    reg node1529_l;
    reg node1530;
    reg node1531;
    reg node1532_r;
    reg node1532_l;
    reg node1533;
    reg node1534;
    reg node1535_r;
    reg node1535_l;
    reg node1536_r;
    reg node1536_l;
    reg node1537_r;
    reg node1537_l;
    reg node1538_r;
    reg node1538_l;
    reg node1539_r;
    reg node1539_l;
    reg node1540;
    reg node1541;
    reg node1542;
    reg node1543;
    reg node1544_r;
    reg node1544_l;
    reg node1545_r;
    reg node1545_l;
    reg node1546;
    reg node1547;
    reg node1548;
    reg node1549_r;
    reg node1549_l;
    reg node1550_r;
    reg node1550_l;
    reg node1551_r;
    reg node1551_l;
    reg node1552_r;
    reg node1552_l;
    reg node1553;
    reg node1554;
    reg node1555;
    reg node1556_r;
    reg node1556_l;
    reg node1557;
    reg node1558_r;
    reg node1558_l;
    reg node1559;
    reg node1560;
    reg node1561_r;
    reg node1561_l;
    reg node1562_r;
    reg node1562_l;
    reg node1563_r;
    reg node1563_l;
    reg node1564;
    reg node1565;
    reg node1566;
    reg node1567_r;
    reg node1567_l;
    reg node1568;
    reg node1569;
    reg node1570_r;
    reg node1570_l;
    reg node1571_r;
    reg node1571_l;
    reg node1572_r;
    reg node1572_l;
    reg node1573_r;
    reg node1573_l;
    reg node1574_r;
    reg node1574_l;
    reg node1575_r;
    reg node1575_l;
    reg node1576;
    reg node1577;
    reg node1578_r;
    reg node1578_l;
    reg node1579;
    reg node1580;
    reg node1581_r;
    reg node1581_l;
    reg node1582_r;
    reg node1582_l;
    reg node1583;
    reg node1584;
    reg node1585_r;
    reg node1585_l;
    reg node1586;
    reg node1587;
    reg node1588_r;
    reg node1588_l;
    reg node1589_r;
    reg node1589_l;
    reg node1590_r;
    reg node1590_l;
    reg node1591;
    reg node1592;
    reg node1593_r;
    reg node1593_l;
    reg node1594;
    reg node1595;
    reg node1596_r;
    reg node1596_l;
    reg node1597_r;
    reg node1597_l;
    reg node1598;
    reg node1599;
    reg node1600_r;
    reg node1600_l;
    reg node1601;
    reg node1602;
    reg node1603_r;
    reg node1603_l;
    reg node1604_r;
    reg node1604_l;
    reg node1605_r;
    reg node1605_l;
    reg node1606_r;
    reg node1606_l;
    reg node1607;
    reg node1608;
    reg node1609_r;
    reg node1609_l;
    reg node1610;
    reg node1611;
    reg node1612_r;
    reg node1612_l;
    reg node1613_r;
    reg node1613_l;
    reg node1614;
    reg node1615;
    reg node1616_r;
    reg node1616_l;
    reg node1617;
    reg node1618;
    reg node1619_r;
    reg node1619_l;
    reg node1620_r;
    reg node1620_l;
    reg node1621_r;
    reg node1621_l;
    reg node1622;
    reg node1623;
    reg node1624_r;
    reg node1624_l;
    reg node1625;
    reg node1626;
    reg node1627_r;
    reg node1627_l;
    reg node1628_r;
    reg node1628_l;
    reg node1629;
    reg node1630;
    reg node1631_r;
    reg node1631_l;
    reg node1632;
    reg node1633;
    reg node1634_r;
    reg node1634_l;
    reg node1635_r;
    reg node1635_l;
    reg node1636_r;
    reg node1636_l;
    reg node1637_r;
    reg node1637_l;
    reg node1638_r;
    reg node1638_l;
    reg node1639;
    reg node1640;
    reg node1641_r;
    reg node1641_l;
    reg node1642;
    reg node1643;
    reg node1644_r;
    reg node1644_l;
    reg node1645;
    reg node1646;
    reg node1647_r;
    reg node1647_l;
    reg node1648_r;
    reg node1648_l;
    reg node1649_r;
    reg node1649_l;
    reg node1650;
    reg node1651;
    reg node1652_r;
    reg node1652_l;
    reg node1653;
    reg node1654;
    reg node1655_r;
    reg node1655_l;
    reg node1656_r;
    reg node1656_l;
    reg node1657;
    reg node1658;
    reg node1659_r;
    reg node1659_l;
    reg node1660;
    reg node1661;
    reg node1662_r;
    reg node1662_l;
    reg node1663_r;
    reg node1663_l;
    reg node1664_r;
    reg node1664_l;
    reg node1665_r;
    reg node1665_l;
    reg node1666;
    reg node1667;
    reg node1668_r;
    reg node1668_l;
    reg node1669;
    reg node1670;
    reg node1671_r;
    reg node1671_l;
    reg node1672_r;
    reg node1672_l;
    reg node1673;
    reg node1674;
    reg node1675_r;
    reg node1675_l;
    reg node1676;
    reg node1677;
    reg node1678_r;
    reg node1678_l;
    reg node1679_r;
    reg node1679_l;
    reg node1680_r;
    reg node1680_l;
    reg node1681;
    reg node1682;
    reg node1683_r;
    reg node1683_l;
    reg node1684;
    reg node1685;
    reg node1686_r;
    reg node1686_l;
    reg node1687_r;
    reg node1687_l;
    reg node1688;
    reg node1689;
    reg node1690_r;
    reg node1690_l;
    reg node1691;
    reg node1692;
    reg result0;
    reg result1;
    reg result2;
    reg result3;
    reg result4;
    reg result5;
    reg result6;
    reg result7;
    reg result8;
    reg result9;

    begin
      node0_r = pixel[406];
      node0_l = ~pixel[406];
      node1_r = node0_l & pixel[414];
      node1_l = node0_l & ~pixel[414];
      node2_r = node1_l & pixel[429];
      node2_l = node1_l & ~pixel[429];
      node3_r = node2_l & pixel[540];
      node3_l = node2_l & ~pixel[540];
      node4_r = node3_l & pixel[260];
      node4_l = node3_l & ~pixel[260];
      node5_r = node4_l & pixel[153];
      node5_l = node4_l & ~pixel[153];
      node6_r = node5_l & pixel[129];
      node6_l = node5_l & ~pixel[129];
      node7_r = node6_l & pixel[464];
      node7_l = node6_l & ~pixel[464];
      node8_r = node7_l & pixel[327];
      node8_l = node7_l & ~pixel[327];
      node9_r = node8_l & pixel[609];
      node9_l = node8_l & ~pixel[609];
      node10 = node9_l;
      node11 = node9_r;
      node12_r = node8_r & pixel[460];
      node12_l = node8_r & ~pixel[460];
      node13 = node12_l;
      node14 = node12_r;
      node15_r = node7_r & pixel[157];
      node15_l = node7_r & ~pixel[157];
      node16_r = node15_l & pixel[267];
      node16_l = node15_l & ~pixel[267];
      node17 = node16_l;
      node18 = node16_r;
      node19_r = node15_r & pixel[654];
      node19_l = node15_r & ~pixel[654];
      node20 = node19_l;
      node21 = node19_r;
      node22_r = node6_r & pixel[217];
      node22_l = node6_r & ~pixel[217];
      node23_r = node22_l & pixel[345];
      node23_l = node22_l & ~pixel[345];
      node24_r = node23_l & pixel[594];
      node24_l = node23_l & ~pixel[594];
      node25 = node24_l;
      node26 = node24_r;
      node27_r = node23_r & pixel[293];
      node27_l = node23_r & ~pixel[293];
      node28 = node27_l;
      node29 = node27_r;
      node30_r = node22_r & pixel[324];
      node30_l = node22_r & ~pixel[324];
      node31_r = node30_l & pixel[512];
      node31_l = node30_l & ~pixel[512];
      node32 = node31_l;
      node33 = node31_r;
      node34_r = node30_r & pixel[467];
      node34_l = node30_r & ~pixel[467];
      node35 = node34_l;
      node36 = node34_r;
      node37_r = node5_r & pixel[267];
      node37_l = node5_r & ~pixel[267];
      node38_r = node37_l & pixel[516];
      node38_l = node37_l & ~pixel[516];
      node39_r = node38_l & pixel[268];
      node39_l = node38_l & ~pixel[268];
      node40_r = node39_l & pixel[319];
      node40_l = node39_l & ~pixel[319];
      node41 = node40_l;
      node42 = node40_r;
      node43_r = node39_r & pixel[295];
      node43_l = node39_r & ~pixel[295];
      node44 = node43_l;
      node45 = node43_r;
      node46_r = node38_r & pixel[459];
      node46_l = node38_r & ~pixel[459];
      node47_r = node46_l & pixel[261];
      node47_l = node46_l & ~pixel[261];
      node48 = node47_l;
      node49 = node47_r;
      node50_r = node46_r & pixel[242];
      node50_l = node46_r & ~pixel[242];
      node51 = node50_l;
      node52 = node50_r;
      node53_r = node37_r & pixel[516];
      node53_l = node37_r & ~pixel[516];
      node54_r = node53_l & pixel[625];
      node54_l = node53_l & ~pixel[625];
      node55_r = node54_l & pixel[351];
      node55_l = node54_l & ~pixel[351];
      node56 = node55_l;
      node57 = node55_r;
      node58_r = node54_r & pixel[329];
      node58_l = node54_r & ~pixel[329];
      node59 = node58_l;
      node60 = node58_r;
      node61_r = node53_r & pixel[376];
      node61_l = node53_r & ~pixel[376];
      node62_r = node61_l & pixel[462];
      node62_l = node61_l & ~pixel[462];
      node63 = node62_l;
      node64 = node62_r;
      node65_r = node61_r & pixel[353];
      node65_l = node61_r & ~pixel[353];
      node66 = node65_l;
      node67 = node65_r;
      node68_r = node4_r & pixel[609];
      node68_l = node4_r & ~pixel[609];
      node69_r = node68_l & pixel[182];
      node69_l = node68_l & ~pixel[182];
      node70_r = node69_l & pixel[483];
      node70_l = node69_l & ~pixel[483];
      node71_r = node70_l & pixel[263];
      node71_l = node70_l & ~pixel[263];
      node72_r = node71_l & pixel[682];
      node72_l = node71_l & ~pixel[682];
      node73 = node72_l;
      node74 = node72_r;
      node75_r = node71_r & pixel[430];
      node75_l = node71_r & ~pixel[430];
      node76 = node75_l;
      node77 = node75_r;
      node78_r = node70_r & pixel[486];
      node78_l = node70_r & ~pixel[486];
      node79_r = node78_l & pixel[371];
      node79_l = node78_l & ~pixel[371];
      node80 = node79_l;
      node81 = node79_r;
      node82_r = node78_r & pixel[528];
      node82_l = node78_r & ~pixel[528];
      node83 = node82_l;
      node84 = node82_r;
      node85_r = node69_r & pixel[634];
      node85_l = node69_r & ~pixel[634];
      node86_r = node85_l & pixel[157];
      node86_l = node85_l & ~pixel[157];
      node87_r = node86_l & pixel[347];
      node87_l = node86_l & ~pixel[347];
      node88 = node87_l;
      node89 = node87_r;
      node90_r = node86_r & pixel[516];
      node90_l = node86_r & ~pixel[516];
      node91 = node90_l;
      node92 = node90_r;
      node93_r = node85_r & pixel[348];
      node93_l = node85_r & ~pixel[348];
      node94_r = node93_l & pixel[571];
      node94_l = node93_l & ~pixel[571];
      node95 = node94_l;
      node96 = node94_r;
      node97_r = node93_r & pixel[551];
      node97_l = node93_r & ~pixel[551];
      node98 = node97_l;
      node99 = node97_r;
      node100_r = node68_r & pixel[542];
      node100_l = node68_r & ~pixel[542];
      node101_r = node100_l & pixel[441];
      node101_l = node100_l & ~pixel[441];
      node102_r = node101_l & pixel[605];
      node102_l = node101_l & ~pixel[605];
      node103_r = node102_l & pixel[255];
      node103_l = node102_l & ~pixel[255];
      node104 = node103_l;
      node105 = node103_r;
      node106_r = node102_r & pixel[369];
      node106_l = node102_r & ~pixel[369];
      node107 = node106_l;
      node108 = node106_r;
      node109_r = node101_r & pixel[267];
      node109_l = node101_r & ~pixel[267];
      node110_r = node109_l & pixel[300];
      node110_l = node109_l & ~pixel[300];
      node111 = node110_l;
      node112 = node110_r;
      node113_r = node109_r & pixel[352];
      node113_l = node109_r & ~pixel[352];
      node114 = node113_l;
      node115 = node113_r;
      node116_r = node100_r & pixel[350];
      node116_l = node100_r & ~pixel[350];
      node117_r = node116_l & pixel[468];
      node117_l = node116_l & ~pixel[468];
      node118_r = node117_l & pixel[599];
      node118_l = node117_l & ~pixel[599];
      node119 = node118_l;
      node120 = node118_r;
      node121_r = node117_r & pixel[487];
      node121_l = node117_r & ~pixel[487];
      node122 = node121_l;
      node123 = node121_r;
      node124_r = node116_r & pixel[430];
      node124_l = node116_r & ~pixel[430];
      node125_r = node124_l & pixel[239];
      node125_l = node124_l & ~pixel[239];
      node126 = node125_l;
      node127 = node125_r;
      node128_r = node124_r & pixel[405];
      node128_l = node124_r & ~pixel[405];
      node129 = node128_l;
      node130 = node128_r;
      node131_r = node3_r & pixel[321];
      node131_l = node3_r & ~pixel[321];
      node132_r = node131_l & pixel[595];
      node132_l = node131_l & ~pixel[595];
      node133_r = node132_l & pixel[482];
      node133_l = node132_l & ~pixel[482];
      node134_r = node133_l & pixel[345];
      node134_l = node133_l & ~pixel[345];
      node135_r = node134_l & pixel[151];
      node135_l = node134_l & ~pixel[151];
      node136_r = node135_l & pixel[158];
      node136_l = node135_l & ~pixel[158];
      node137 = node136_l;
      node138 = node136_r;
      node139_r = node135_r & pixel[400];
      node139_l = node135_r & ~pixel[400];
      node140 = node139_l;
      node141 = node139_r;
      node142_r = node134_r & pixel[374];
      node142_l = node134_r & ~pixel[374];
      node143_r = node142_l & pixel[483];
      node143_l = node142_l & ~pixel[483];
      node144 = node143_l;
      node145 = node143_r;
      node146_r = node142_r & pixel[436];
      node146_l = node142_r & ~pixel[436];
      node147 = node146_l;
      node148 = node146_r;
      node149_r = node133_r & pixel[155];
      node149_l = node133_r & ~pixel[155];
      node150_r = node149_l & pixel[185];
      node150_l = node149_l & ~pixel[185];
      node151_r = node150_l & pixel[410];
      node151_l = node150_l & ~pixel[410];
      node152 = node151_l;
      node153 = node151_r;
      node154_r = node150_r & pixel[352];
      node154_l = node150_r & ~pixel[352];
      node155 = node154_l;
      node156 = node154_r;
      node157_r = node149_r & pixel[444];
      node157_l = node149_r & ~pixel[444];
      node158_r = node157_l & pixel[524];
      node158_l = node157_l & ~pixel[524];
      node159 = node158_l;
      node160 = node158_r;
      node161_r = node157_r & pixel[274];
      node161_l = node157_r & ~pixel[274];
      node162 = node161_l;
      node163 = node161_r;
      node164_r = node132_r & pixel[490];
      node164_l = node132_r & ~pixel[490];
      node165_r = node164_l & pixel[290];
      node165_l = node164_l & ~pixel[290];
      node166_r = node165_l & pixel[416];
      node166_l = node165_l & ~pixel[416];
      node167_r = node166_l & pixel[484];
      node167_l = node166_l & ~pixel[484];
      node168 = node167_l;
      node169 = node167_r;
      node170 = node166_r;
      node171_r = node165_r & pixel[370];
      node171_l = node165_r & ~pixel[370];
      node172_r = node171_l & pixel[684];
      node172_l = node171_l & ~pixel[684];
      node173 = node172_l;
      node174 = node172_r;
      node175_r = node171_r & pixel[513];
      node175_l = node171_r & ~pixel[513];
      node176 = node175_l;
      node177 = node175_r;
      node178_r = node164_r & pixel[680];
      node178_l = node164_r & ~pixel[680];
      node179_r = node178_l & pixel[398];
      node179_l = node178_l & ~pixel[398];
      node180_r = node179_l & pixel[684];
      node180_l = node179_l & ~pixel[684];
      node181 = node180_l;
      node182 = node180_r;
      node183_r = node179_r & pixel[300];
      node183_l = node179_r & ~pixel[300];
      node184 = node183_l;
      node185 = node183_r;
      node186_r = node178_r & pixel[634];
      node186_l = node178_r & ~pixel[634];
      node187_r = node186_l & pixel[180];
      node187_l = node186_l & ~pixel[180];
      node188 = node187_l;
      node189 = node187_r;
      node190_r = node186_r & pixel[598];
      node190_l = node186_r & ~pixel[598];
      node191 = node190_l;
      node192 = node190_r;
      node193_r = node131_r & pixel[179];
      node193_l = node131_r & ~pixel[179];
      node194_r = node193_l & pixel[403];
      node194_l = node193_l & ~pixel[403];
      node195_r = node194_l & pixel[301];
      node195_l = node194_l & ~pixel[301];
      node196_r = node195_l & pixel[151];
      node196_l = node195_l & ~pixel[151];
      node197_r = node196_l & pixel[351];
      node197_l = node196_l & ~pixel[351];
      node198 = node197_l;
      node199 = node197_r;
      node200_r = node196_r & pixel[480];
      node200_l = node196_r & ~pixel[480];
      node201 = node200_l;
      node202 = node200_r;
      node203_r = node195_r & pixel[464];
      node203_l = node195_r & ~pixel[464];
      node204_r = node203_l & pixel[470];
      node204_l = node203_l & ~pixel[470];
      node205 = node204_l;
      node206 = node204_r;
      node207_r = node203_r & pixel[371];
      node207_l = node203_r & ~pixel[371];
      node208 = node207_l;
      node209 = node207_r;
      node210_r = node194_r & pixel[245];
      node210_l = node194_r & ~pixel[245];
      node211_r = node210_l & pixel[127];
      node211_l = node210_l & ~pixel[127];
      node212_r = node211_l & pixel[431];
      node212_l = node211_l & ~pixel[431];
      node213 = node212_l;
      node214 = node212_r;
      node215_r = node211_r & pixel[351];
      node215_l = node211_r & ~pixel[351];
      node216 = node215_l;
      node217 = node215_r;
      node218_r = node210_r & pixel[495];
      node218_l = node210_r & ~pixel[495];
      node219_r = node218_l & pixel[355];
      node219_l = node218_l & ~pixel[355];
      node220 = node219_l;
      node221 = node219_r;
      node222_r = node218_r & pixel[247];
      node222_l = node218_r & ~pixel[247];
      node223 = node222_l;
      node224 = node222_r;
      node225_r = node193_r & pixel[270];
      node225_l = node193_r & ~pixel[270];
      node226_r = node225_l & pixel[158];
      node226_l = node225_l & ~pixel[158];
      node227_r = node226_l & pixel[432];
      node227_l = node226_l & ~pixel[432];
      node228_r = node227_l & pixel[637];
      node228_l = node227_l & ~pixel[637];
      node229 = node228_l;
      node230 = node228_r;
      node231_r = node227_r & pixel[439];
      node231_l = node227_r & ~pixel[439];
      node232 = node231_l;
      node233 = node231_r;
      node234_r = node226_r & pixel[240];
      node234_l = node226_r & ~pixel[240];
      node235_r = node234_l & pixel[361];
      node235_l = node234_l & ~pixel[361];
      node236 = node235_l;
      node237 = node235_r;
      node238_r = node234_r & pixel[215];
      node238_l = node234_r & ~pixel[215];
      node239 = node238_l;
      node240 = node238_r;
      node241_r = node225_r & pixel[631];
      node241_l = node225_r & ~pixel[631];
      node242_r = node241_l & pixel[525];
      node242_l = node241_l & ~pixel[525];
      node243_r = node242_l & pixel[486];
      node243_l = node242_l & ~pixel[486];
      node244 = node243_l;
      node245 = node243_r;
      node246_r = node242_r & pixel[519];
      node246_l = node242_r & ~pixel[519];
      node247 = node246_l;
      node248 = node246_r;
      node249_r = node241_r & pixel[295];
      node249_l = node241_r & ~pixel[295];
      node250_r = node249_l & pixel[126];
      node250_l = node249_l & ~pixel[126];
      node251 = node250_l;
      node252 = node250_r;
      node253_r = node249_r & pixel[162];
      node253_l = node249_r & ~pixel[162];
      node254 = node253_l;
      node255 = node253_r;
      node256_r = node2_r & pixel[655];
      node256_l = node2_r & ~pixel[655];
      node257_r = node256_l & pixel[325];
      node257_l = node256_l & ~pixel[325];
      node258_r = node257_l & pixel[130];
      node258_l = node257_l & ~pixel[130];
      node259_r = node258_l & pixel[355];
      node259_l = node258_l & ~pixel[355];
      node260_r = node259_l & pixel[247];
      node260_l = node259_l & ~pixel[247];
      node261_r = node260_l & pixel[99];
      node261_l = node260_l & ~pixel[99];
      node262_r = node261_l & pixel[542];
      node262_l = node261_l & ~pixel[542];
      node263 = node262_l;
      node264 = node262_r;
      node265_r = node261_r & pixel[213];
      node265_l = node261_r & ~pixel[213];
      node266 = node265_l;
      node267 = node265_r;
      node268_r = node260_r & pixel[678];
      node268_l = node260_r & ~pixel[678];
      node269_r = node268_l & pixel[356];
      node269_l = node268_l & ~pixel[356];
      node270 = node269_l;
      node271 = node269_r;
      node272 = node268_r;
      node273_r = node259_r & pixel[213];
      node273_l = node259_r & ~pixel[213];
      node274_r = node273_l & pixel[570];
      node274_l = node273_l & ~pixel[570];
      node275_r = node274_l & pixel[712];
      node275_l = node274_l & ~pixel[712];
      node276 = node275_l;
      node277 = node275_r;
      node278_r = node274_r & pixel[237];
      node278_l = node274_r & ~pixel[237];
      node279 = node278_l;
      node280 = node278_r;
      node281_r = node273_r & pixel[461];
      node281_l = node273_r & ~pixel[461];
      node282_r = node281_l & pixel[384];
      node282_l = node281_l & ~pixel[384];
      node283 = node282_l;
      node284 = node282_r;
      node285_r = node281_r & pixel[537];
      node285_l = node281_r & ~pixel[537];
      node286 = node285_l;
      node287 = node285_r;
      node288_r = node258_r & pixel[592];
      node288_l = node258_r & ~pixel[592];
      node289_r = node288_l & pixel[215];
      node289_l = node288_l & ~pixel[215];
      node290_r = node289_l & pixel[125];
      node290_l = node289_l & ~pixel[125];
      node291_r = node290_l & pixel[357];
      node291_l = node290_l & ~pixel[357];
      node292 = node291_l;
      node293 = node291_r;
      node294_r = node290_r & pixel[538];
      node294_l = node290_r & ~pixel[538];
      node295 = node294_l;
      node296 = node294_r;
      node297_r = node289_r & pixel[565];
      node297_l = node289_r & ~pixel[565];
      node298_r = node297_l & pixel[517];
      node298_l = node297_l & ~pixel[517];
      node299 = node298_l;
      node300 = node298_r;
      node301_r = node297_r & pixel[105];
      node301_l = node297_r & ~pixel[105];
      node302 = node301_l;
      node303 = node301_r;
      node304_r = node288_r & pixel[378];
      node304_l = node288_r & ~pixel[378];
      node305_r = node304_l & pixel[459];
      node305_l = node304_l & ~pixel[459];
      node306_r = node305_l & pixel[291];
      node306_l = node305_l & ~pixel[291];
      node307 = node306_l;
      node308 = node306_r;
      node309 = node305_r;
      node310 = node304_r;
      node311_r = node257_r & pixel[462];
      node311_l = node257_r & ~pixel[462];
      node312_r = node311_l & pixel[718];
      node312_l = node311_l & ~pixel[718];
      node313_r = node312_l & pixel[599];
      node313_l = node312_l & ~pixel[599];
      node314_r = node313_l & pixel[515];
      node314_l = node313_l & ~pixel[515];
      node315_r = node314_l & pixel[268];
      node315_l = node314_l & ~pixel[268];
      node316 = node315_l;
      node317 = node315_r;
      node318_r = node314_r & pixel[716];
      node318_l = node314_r & ~pixel[716];
      node319 = node318_l;
      node320 = node318_r;
      node321_r = node313_r & pixel[351];
      node321_l = node313_r & ~pixel[351];
      node322_r = node321_l & pixel[628];
      node322_l = node321_l & ~pixel[628];
      node323 = node322_l;
      node324 = node322_r;
      node325_r = node321_r & pixel[567];
      node325_l = node321_r & ~pixel[567];
      node326 = node325_l;
      node327 = node325_r;
      node328_r = node312_r & pixel[264];
      node328_l = node312_r & ~pixel[264];
      node329_r = node328_l & pixel[374];
      node329_l = node328_l & ~pixel[374];
      node330 = node329_l;
      node331_r = node329_r & pixel[233];
      node331_l = node329_r & ~pixel[233];
      node332 = node331_l;
      node333 = node331_r;
      node334_r = node328_r & pixel[233];
      node334_l = node328_r & ~pixel[233];
      node335_r = node334_l & pixel[690];
      node335_l = node334_l & ~pixel[690];
      node336 = node335_l;
      node337 = node335_r;
      node338_r = node334_r & pixel[369];
      node338_l = node334_r & ~pixel[369];
      node339 = node338_l;
      node340 = node338_r;
      node341_r = node311_r & pixel[99];
      node341_l = node311_r & ~pixel[99];
      node342_r = node341_l & pixel[161];
      node342_l = node341_l & ~pixel[161];
      node343_r = node342_l & pixel[720];
      node343_l = node342_l & ~pixel[720];
      node344_r = node343_l & pixel[373];
      node344_l = node343_l & ~pixel[373];
      node345 = node344_l;
      node346 = node344_r;
      node347_r = node343_r & pixel[629];
      node347_l = node343_r & ~pixel[629];
      node348 = node347_l;
      node349 = node347_r;
      node350_r = node342_r & pixel[212];
      node350_l = node342_r & ~pixel[212];
      node351_r = node350_l & pixel[623];
      node351_l = node350_l & ~pixel[623];
      node352 = node351_l;
      node353 = node351_r;
      node354_r = node350_r & pixel[467];
      node354_l = node350_r & ~pixel[467];
      node355 = node354_l;
      node356 = node354_r;
      node357_r = node341_r & pixel[344];
      node357_l = node341_r & ~pixel[344];
      node358_r = node357_l & pixel[291];
      node358_l = node357_l & ~pixel[291];
      node359_r = node358_l & pixel[398];
      node359_l = node358_l & ~pixel[398];
      node360 = node359_l;
      node361 = node359_r;
      node362_r = node358_r & pixel[539];
      node362_l = node358_r & ~pixel[539];
      node363 = node362_l;
      node364 = node362_r;
      node365_r = node357_r & pixel[156];
      node365_l = node357_r & ~pixel[156];
      node366 = node365_l;
      node367_r = node365_r & pixel[289];
      node367_l = node365_r & ~pixel[289];
      node368 = node367_l;
      node369 = node367_r;
      node370_r = node256_r & pixel[440];
      node370_l = node256_r & ~pixel[440];
      node371_r = node370_l & pixel[411];
      node371_l = node370_l & ~pixel[411];
      node372_r = node371_l & pixel[409];
      node372_l = node371_l & ~pixel[409];
      node373_r = node372_l & pixel[237];
      node373_l = node372_l & ~pixel[237];
      node374_r = node373_l & pixel[578];
      node374_l = node373_l & ~pixel[578];
      node375_r = node374_l & pixel[220];
      node375_l = node374_l & ~pixel[220];
      node376 = node375_l;
      node377 = node375_r;
      node378_r = node374_r & pixel[153];
      node378_l = node374_r & ~pixel[153];
      node379 = node378_l;
      node380 = node378_r;
      node381_r = node373_r & pixel[131];
      node381_l = node373_r & ~pixel[131];
      node382_r = node381_l & pixel[500];
      node382_l = node381_l & ~pixel[500];
      node383 = node382_l;
      node384 = node382_r;
      node385_r = node381_r & pixel[207];
      node385_l = node381_r & ~pixel[207];
      node386 = node385_l;
      node387 = node385_r;
      node388_r = node372_r & pixel[545];
      node388_l = node372_r & ~pixel[545];
      node389_r = node388_l & pixel[298];
      node389_l = node388_l & ~pixel[298];
      node390_r = node389_l & pixel[269];
      node390_l = node389_l & ~pixel[269];
      node391 = node390_l;
      node392 = node390_r;
      node393_r = node389_r & pixel[542];
      node393_l = node389_r & ~pixel[542];
      node394 = node393_l;
      node395 = node393_r;
      node396_r = node388_r & pixel[126];
      node396_l = node388_r & ~pixel[126];
      node397_r = node396_l & pixel[296];
      node397_l = node396_l & ~pixel[296];
      node398 = node397_l;
      node399 = node397_r;
      node400_r = node396_r & pixel[602];
      node400_l = node396_r & ~pixel[602];
      node401 = node400_l;
      node402 = node400_r;
      node403_r = node371_r & pixel[158];
      node403_l = node371_r & ~pixel[158];
      node404_r = node403_l & pixel[460];
      node404_l = node403_l & ~pixel[460];
      node405_r = node404_l & pixel[300];
      node405_l = node404_l & ~pixel[300];
      node406_r = node405_l & pixel[350];
      node406_l = node405_l & ~pixel[350];
      node407 = node406_l;
      node408 = node406_r;
      node409_r = node405_r & pixel[624];
      node409_l = node405_r & ~pixel[624];
      node410 = node409_l;
      node411 = node409_r;
      node412_r = node404_r & pixel[212];
      node412_l = node404_r & ~pixel[212];
      node413_r = node412_l & pixel[582];
      node413_l = node412_l & ~pixel[582];
      node414 = node413_l;
      node415 = node413_r;
      node416_r = node412_r & pixel[596];
      node416_l = node412_r & ~pixel[596];
      node417 = node416_l;
      node418 = node416_r;
      node419_r = node403_r & pixel[152];
      node419_l = node403_r & ~pixel[152];
      node420_r = node419_l & pixel[303];
      node420_l = node419_l & ~pixel[303];
      node421_r = node420_l & pixel[551];
      node421_l = node420_l & ~pixel[551];
      node422 = node421_l;
      node423 = node421_r;
      node424_r = node420_r & pixel[428];
      node424_l = node420_r & ~pixel[428];
      node425 = node424_l;
      node426 = node424_r;
      node427_r = node419_r & pixel[402];
      node427_l = node419_r & ~pixel[402];
      node428_r = node427_l & pixel[379];
      node428_l = node427_l & ~pixel[379];
      node429 = node428_l;
      node430 = node428_r;
      node431_r = node427_r & pixel[464];
      node431_l = node427_r & ~pixel[464];
      node432 = node431_l;
      node433 = node431_r;
      node434_r = node370_r & pixel[381];
      node434_l = node370_r & ~pixel[381];
      node435_r = node434_l & pixel[484];
      node435_l = node434_l & ~pixel[484];
      node436_r = node435_l & pixel[205];
      node436_l = node435_l & ~pixel[205];
      node437_r = node436_l & pixel[545];
      node437_l = node436_l & ~pixel[545];
      node438_r = node437_l & pixel[242];
      node438_l = node437_l & ~pixel[242];
      node439 = node438_l;
      node440 = node438_r;
      node441_r = node437_r & pixel[460];
      node441_l = node437_r & ~pixel[460];
      node442 = node441_l;
      node443 = node441_r;
      node444_r = node436_r & pixel[515];
      node444_l = node436_r & ~pixel[515];
      node445_r = node444_l & pixel[348];
      node445_l = node444_l & ~pixel[348];
      node446 = node445_l;
      node447 = node445_r;
      node448_r = node444_r & pixel[274];
      node448_l = node444_r & ~pixel[274];
      node449 = node448_l;
      node450 = node448_r;
      node451_r = node435_r & pixel[401];
      node451_l = node435_r & ~pixel[401];
      node452_r = node451_l & pixel[626];
      node452_l = node451_l & ~pixel[626];
      node453_r = node452_l & pixel[573];
      node453_l = node452_l & ~pixel[573];
      node454 = node453_l;
      node455 = node453_r;
      node456_r = node452_r & pixel[377];
      node456_l = node452_r & ~pixel[377];
      node457 = node456_l;
      node458 = node456_r;
      node459_r = node451_r & pixel[443];
      node459_l = node451_r & ~pixel[443];
      node460_r = node459_l & pixel[709];
      node460_l = node459_l & ~pixel[709];
      node461 = node460_l;
      node462 = node460_r;
      node463 = node459_r;
      node464_r = node434_r & pixel[327];
      node464_l = node434_r & ~pixel[327];
      node465_r = node464_l & pixel[290];
      node465_l = node464_l & ~pixel[290];
      node466_r = node465_l & pixel[343];
      node466_l = node465_l & ~pixel[343];
      node467_r = node466_l & pixel[717];
      node467_l = node466_l & ~pixel[717];
      node468 = node467_l;
      node469 = node467_r;
      node470_r = node466_r & pixel[412];
      node470_l = node466_r & ~pixel[412];
      node471 = node470_l;
      node472 = node470_r;
      node473_r = node465_r & pixel[486];
      node473_l = node465_r & ~pixel[486];
      node474_r = node473_l & pixel[259];
      node474_l = node473_l & ~pixel[259];
      node475 = node474_l;
      node476 = node474_r;
      node477_r = node473_r & pixel[578];
      node477_l = node473_r & ~pixel[578];
      node478 = node477_l;
      node479 = node477_r;
      node480_r = node464_r & pixel[183];
      node480_l = node464_r & ~pixel[183];
      node481_r = node480_l & pixel[622];
      node481_l = node480_l & ~pixel[622];
      node482_r = node481_l & pixel[266];
      node482_l = node481_l & ~pixel[266];
      node483 = node482_l;
      node484 = node482_r;
      node485 = node481_r;
      node486_r = node480_r & pixel[549];
      node486_l = node480_r & ~pixel[549];
      node487_r = node486_l & pixel[497];
      node487_l = node486_l & ~pixel[497];
      node488 = node487_l;
      node489 = node487_r;
      node490_r = node486_r & pixel[489];
      node490_l = node486_r & ~pixel[489];
      node491 = node490_l;
      node492 = node490_r;
      node493_r = node1_r & pixel[490];
      node493_l = node1_r & ~pixel[490];
      node494_r = node493_l & pixel[245];
      node494_l = node493_l & ~pixel[245];
      node495_r = node494_l & pixel[352];
      node495_l = node494_l & ~pixel[352];
      node496_r = node495_l & pixel[436];
      node496_l = node495_l & ~pixel[436];
      node497_r = node496_l & pixel[598];
      node497_l = node496_l & ~pixel[598];
      node498_r = node497_l & pixel[511];
      node498_l = node497_l & ~pixel[511];
      node499_r = node498_l & pixel[542];
      node499_l = node498_l & ~pixel[542];
      node500_r = node499_l & pixel[510];
      node500_l = node499_l & ~pixel[510];
      node501 = node500_l;
      node502 = node500_r;
      node503_r = node499_r & pixel[300];
      node503_l = node499_r & ~pixel[300];
      node504 = node503_l;
      node505 = node503_r;
      node506_r = node498_r & pixel[351];
      node506_l = node498_r & ~pixel[351];
      node507_r = node506_l & pixel[742];
      node507_l = node506_l & ~pixel[742];
      node508 = node507_l;
      node509 = node507_r;
      node510 = node506_r;
      node511_r = node497_r & pixel[656];
      node511_l = node497_r & ~pixel[656];
      node512_r = node511_l & pixel[214];
      node512_l = node511_l & ~pixel[214];
      node513_r = node512_l & pixel[69];
      node513_l = node512_l & ~pixel[69];
      node514 = node513_l;
      node515 = node513_r;
      node516_r = node512_r & pixel[128];
      node516_l = node512_r & ~pixel[128];
      node517 = node516_l;
      node518 = node516_r;
      node519_r = node511_r & pixel[545];
      node519_l = node511_r & ~pixel[545];
      node520_r = node519_l & pixel[295];
      node520_l = node519_l & ~pixel[295];
      node521 = node520_l;
      node522 = node520_r;
      node523_r = node519_r & pixel[552];
      node523_l = node519_r & ~pixel[552];
      node524 = node523_l;
      node525 = node523_r;
      node526_r = node496_r & pixel[372];
      node526_l = node496_r & ~pixel[372];
      node527_r = node526_l & pixel[325];
      node527_l = node526_l & ~pixel[325];
      node528_r = node527_l & pixel[494];
      node528_l = node527_l & ~pixel[494];
      node529_r = node528_l & pixel[539];
      node529_l = node528_l & ~pixel[539];
      node530 = node529_l;
      node531 = node529_r;
      node532_r = node528_r & pixel[75];
      node532_l = node528_r & ~pixel[75];
      node533 = node532_l;
      node534 = node532_r;
      node535_r = node527_r & pixel[456];
      node535_l = node527_r & ~pixel[456];
      node536 = node535_l;
      node537 = node535_r;
      node538_r = node526_r & pixel[243];
      node538_l = node526_r & ~pixel[243];
      node539_r = node538_l & pixel[432];
      node539_l = node538_l & ~pixel[432];
      node540 = node539_l;
      node541_r = node539_r & pixel[608];
      node541_l = node539_r & ~pixel[608];
      node542 = node541_l;
      node543 = node541_r;
      node544 = node538_r;
      node545_r = node495_r & pixel[212];
      node545_l = node495_r & ~pixel[212];
      node546_r = node545_l & pixel[153];
      node546_l = node545_l & ~pixel[153];
      node547_r = node546_l & pixel[458];
      node547_l = node546_l & ~pixel[458];
      node548_r = node547_l & pixel[466];
      node548_l = node547_l & ~pixel[466];
      node549_r = node548_l & pixel[239];
      node549_l = node548_l & ~pixel[239];
      node550 = node549_l;
      node551 = node549_r;
      node552_r = node548_r & pixel[624];
      node552_l = node548_r & ~pixel[624];
      node553 = node552_l;
      node554 = node552_r;
      node555_r = node547_r & pixel[688];
      node555_l = node547_r & ~pixel[688];
      node556 = node555_l;
      node557_r = node555_r & pixel[292];
      node557_l = node555_r & ~pixel[292];
      node558 = node557_l;
      node559 = node557_r;
      node560_r = node546_r & pixel[238];
      node560_l = node546_r & ~pixel[238];
      node561_r = node560_l & pixel[348];
      node561_l = node560_l & ~pixel[348];
      node562_r = node561_l & pixel[578];
      node562_l = node561_l & ~pixel[578];
      node563 = node562_l;
      node564 = node562_r;
      node565_r = node561_r & pixel[628];
      node565_l = node561_r & ~pixel[628];
      node566 = node565_l;
      node567 = node565_r;
      node568_r = node560_r & pixel[546];
      node568_l = node560_r & ~pixel[546];
      node569_r = node568_l & pixel[265];
      node569_l = node568_l & ~pixel[265];
      node570 = node569_l;
      node571 = node569_r;
      node572 = node568_r;
      node573_r = node545_r & pixel[235];
      node573_l = node545_r & ~pixel[235];
      node574_r = node573_l & pixel[261];
      node574_l = node573_l & ~pixel[261];
      node575_r = node574_l & pixel[638];
      node575_l = node574_l & ~pixel[638];
      node576_r = node575_l & pixel[104];
      node576_l = node575_l & ~pixel[104];
      node577 = node576_l;
      node578 = node576_r;
      node579_r = node575_r & pixel[579];
      node579_l = node575_r & ~pixel[579];
      node580 = node579_l;
      node581 = node579_r;
      node582_r = node574_r & pixel[269];
      node582_l = node574_r & ~pixel[269];
      node583_r = node582_l & pixel[186];
      node583_l = node582_l & ~pixel[186];
      node584 = node583_l;
      node585 = node583_r;
      node586_r = node582_r & pixel[348];
      node586_l = node582_r & ~pixel[348];
      node587 = node586_l;
      node588 = node586_r;
      node589_r = node573_r & pixel[347];
      node589_l = node573_r & ~pixel[347];
      node590_r = node589_l & pixel[348];
      node590_l = node589_l & ~pixel[348];
      node591_r = node590_l & pixel[480];
      node591_l = node590_l & ~pixel[480];
      node592 = node591_l;
      node593 = node591_r;
      node594_r = node590_r & pixel[402];
      node594_l = node590_r & ~pixel[402];
      node595 = node594_l;
      node596 = node594_r;
      node597_r = node589_r & pixel[495];
      node597_l = node589_r & ~pixel[495];
      node598_r = node597_l & pixel[244];
      node598_l = node597_l & ~pixel[244];
      node599 = node598_l;
      node600 = node598_r;
      node601_r = node597_r & pixel[272];
      node601_l = node597_r & ~pixel[272];
      node602 = node601_l;
      node603 = node601_r;
      node604_r = node494_r & pixel[712];
      node604_l = node494_r & ~pixel[712];
      node605_r = node604_l & pixel[482];
      node605_l = node604_l & ~pixel[482];
      node606_r = node605_l & pixel[456];
      node606_l = node605_l & ~pixel[456];
      node607_r = node606_l & pixel[355];
      node607_l = node606_l & ~pixel[355];
      node608_r = node607_l & pixel[555];
      node608_l = node607_l & ~pixel[555];
      node609_r = node608_l & pixel[525];
      node609_l = node608_l & ~pixel[525];
      node610 = node609_l;
      node611 = node609_r;
      node612 = node608_r;
      node613_r = node607_r & pixel[269];
      node613_l = node607_r & ~pixel[269];
      node614_r = node613_l & pixel[624];
      node614_l = node613_l & ~pixel[624];
      node615 = node614_l;
      node616 = node614_r;
      node617_r = node613_r & pixel[188];
      node617_l = node613_r & ~pixel[188];
      node618 = node617_l;
      node619 = node617_r;
      node620_r = node606_r & pixel[555];
      node620_l = node606_r & ~pixel[555];
      node621_r = node620_l & pixel[228];
      node621_l = node620_l & ~pixel[228];
      node622 = node621_l;
      node623_r = node621_r & pixel[685];
      node623_l = node621_r & ~pixel[685];
      node624 = node623_l;
      node625 = node623_r;
      node626_r = node620_r & pixel[399];
      node626_l = node620_r & ~pixel[399];
      node627 = node626_l;
      node628 = node626_r;
      node629_r = node605_r & pixel[434];
      node629_l = node605_r & ~pixel[434];
      node630_r = node629_l & pixel[386];
      node630_l = node629_l & ~pixel[386];
      node631_r = node630_l & pixel[323];
      node631_l = node630_l & ~pixel[323];
      node632_r = node631_l & pixel[328];
      node632_l = node631_l & ~pixel[328];
      node633 = node632_l;
      node634 = node632_r;
      node635_r = node631_r & pixel[541];
      node635_l = node631_r & ~pixel[541];
      node636 = node635_l;
      node637 = node635_r;
      node638_r = node630_r & pixel[311];
      node638_l = node630_r & ~pixel[311];
      node639_r = node638_l & pixel[379];
      node639_l = node638_l & ~pixel[379];
      node640 = node639_l;
      node641 = node639_r;
      node642_r = node638_r & pixel[400];
      node642_l = node638_r & ~pixel[400];
      node643 = node642_l;
      node644 = node642_r;
      node645_r = node629_r & pixel[459];
      node645_l = node629_r & ~pixel[459];
      node646 = node645_l;
      node647_r = node645_r & pixel[291];
      node647_l = node645_r & ~pixel[291];
      node648 = node647_l;
      node649 = node647_r;
      node650_r = node604_r & pixel[183];
      node650_l = node604_r & ~pixel[183];
      node651 = node650_l;
      node652_r = node650_r & pixel[353];
      node652_l = node650_r & ~pixel[353];
      node653_r = node652_l & pixel[575];
      node653_l = node652_l & ~pixel[575];
      node654 = node653_l;
      node655_r = node653_r & pixel[574];
      node655_l = node653_r & ~pixel[574];
      node656 = node655_l;
      node657 = node655_r;
      node658_r = node652_r & pixel[411];
      node658_l = node652_r & ~pixel[411];
      node659 = node658_l;
      node660_r = node658_r & pixel[202];
      node660_l = node658_r & ~pixel[202];
      node661 = node660_l;
      node662 = node660_r;
      node663_r = node493_r & pixel[436];
      node663_l = node493_r & ~pixel[436];
      node664_r = node663_l & pixel[371];
      node664_l = node663_l & ~pixel[371];
      node665_r = node664_l & pixel[376];
      node665_l = node664_l & ~pixel[376];
      node666_r = node665_l & pixel[695];
      node666_l = node665_l & ~pixel[695];
      node667_r = node666_l & pixel[707];
      node667_l = node666_l & ~pixel[707];
      node668_r = node667_l & pixel[551];
      node668_l = node667_l & ~pixel[551];
      node669_r = node668_l & pixel[272];
      node669_l = node668_l & ~pixel[272];
      node670 = node669_l;
      node671 = node669_r;
      node672_r = node668_r & pixel[156];
      node672_l = node668_r & ~pixel[156];
      node673 = node672_l;
      node674 = node672_r;
      node675 = node667_r;
      node676 = node666_r;
      node677_r = node665_r & pixel[302];
      node677_l = node665_r & ~pixel[302];
      node678_r = node677_l & pixel[287];
      node678_l = node677_l & ~pixel[287];
      node679_r = node678_l & pixel[301];
      node679_l = node678_l & ~pixel[301];
      node680_r = node679_l & pixel[319];
      node680_l = node679_l & ~pixel[319];
      node681 = node680_l;
      node682 = node680_r;
      node683 = node679_r;
      node684 = node678_r;
      node685_r = node677_r & pixel[261];
      node685_l = node677_r & ~pixel[261];
      node686 = node685_l;
      node687 = node685_r;
      node688_r = node664_r & pixel[538];
      node688_l = node664_r & ~pixel[538];
      node689_r = node688_l & pixel[425];
      node689_l = node688_l & ~pixel[425];
      node690_r = node689_l & pixel[527];
      node690_l = node689_l & ~pixel[527];
      node691_r = node690_l & pixel[544];
      node691_l = node690_l & ~pixel[544];
      node692_r = node691_l & pixel[268];
      node692_l = node691_l & ~pixel[268];
      node693 = node692_l;
      node694 = node692_r;
      node695_r = node691_r & pixel[553];
      node695_l = node691_r & ~pixel[553];
      node696 = node695_l;
      node697 = node695_r;
      node698_r = node690_r & pixel[319];
      node698_l = node690_r & ~pixel[319];
      node699 = node698_l;
      node700_r = node698_r & pixel[239];
      node700_l = node698_r & ~pixel[239];
      node701 = node700_l;
      node702 = node700_r;
      node703_r = node689_r & pixel[525];
      node703_l = node689_r & ~pixel[525];
      node704_r = node703_l & pixel[411];
      node704_l = node703_l & ~pixel[411];
      node705 = node704_l;
      node706 = node704_r;
      node707_r = node703_r & pixel[240];
      node707_l = node703_r & ~pixel[240];
      node708 = node707_l;
      node709 = node707_r;
      node710_r = node688_r & pixel[186];
      node710_l = node688_r & ~pixel[186];
      node711_r = node710_l & pixel[241];
      node711_l = node710_l & ~pixel[241];
      node712_r = node711_l & pixel[231];
      node712_l = node711_l & ~pixel[231];
      node713_r = node712_l & pixel[581];
      node713_l = node712_l & ~pixel[581];
      node714 = node713_l;
      node715 = node713_r;
      node716 = node712_r;
      node717_r = node711_r & pixel[409];
      node717_l = node711_r & ~pixel[409];
      node718 = node717_l;
      node719_r = node717_r & pixel[230];
      node719_l = node717_r & ~pixel[230];
      node720 = node719_l;
      node721 = node719_r;
      node722_r = node710_r & pixel[427];
      node722_l = node710_r & ~pixel[427];
      node723_r = node722_l & pixel[188];
      node723_l = node722_l & ~pixel[188];
      node724 = node723_l;
      node725 = node723_r;
      node726_r = node722_r & pixel[611];
      node726_l = node722_r & ~pixel[611];
      node727_r = node726_l & pixel[569];
      node727_l = node726_l & ~pixel[569];
      node728 = node727_l;
      node729 = node727_r;
      node730 = node726_r;
      node731_r = node663_r & pixel[299];
      node731_l = node663_r & ~pixel[299];
      node732_r = node731_l & pixel[621];
      node732_l = node731_l & ~pixel[621];
      node733_r = node732_l & pixel[296];
      node733_l = node732_l & ~pixel[296];
      node734_r = node733_l & pixel[303];
      node734_l = node733_l & ~pixel[303];
      node735_r = node734_l & pixel[272];
      node735_l = node734_l & ~pixel[272];
      node736_r = node735_l & pixel[549];
      node736_l = node735_l & ~pixel[549];
      node737 = node736_l;
      node738 = node736_r;
      node739_r = node735_r & pixel[469];
      node739_l = node735_r & ~pixel[469];
      node740 = node739_l;
      node741 = node739_r;
      node742_r = node734_r & pixel[347];
      node742_l = node734_r & ~pixel[347];
      node743_r = node742_l & pixel[342];
      node743_l = node742_l & ~pixel[342];
      node744 = node743_l;
      node745 = node743_r;
      node746_r = node742_r & pixel[388];
      node746_l = node742_r & ~pixel[388];
      node747 = node746_l;
      node748 = node746_r;
      node749_r = node733_r & pixel[572];
      node749_l = node733_r & ~pixel[572];
      node750_r = node749_l & pixel[286];
      node750_l = node749_l & ~pixel[286];
      node751_r = node750_l & pixel[204];
      node751_l = node750_l & ~pixel[204];
      node752 = node751_l;
      node753 = node751_r;
      node754_r = node750_r & pixel[636];
      node754_l = node750_r & ~pixel[636];
      node755 = node754_l;
      node756 = node754_r;
      node757_r = node749_r & pixel[386];
      node757_l = node749_r & ~pixel[386];
      node758_r = node757_l & pixel[627];
      node758_l = node757_l & ~pixel[627];
      node759 = node758_l;
      node760 = node758_r;
      node761_r = node757_r & pixel[330];
      node761_l = node757_r & ~pixel[330];
      node762 = node761_l;
      node763 = node761_r;
      node764_r = node732_r & pixel[400];
      node764_l = node732_r & ~pixel[400];
      node765_r = node764_l & pixel[261];
      node765_l = node764_l & ~pixel[261];
      node766_r = node765_l & pixel[276];
      node766_l = node765_l & ~pixel[276];
      node767_r = node766_l & pixel[208];
      node767_l = node766_l & ~pixel[208];
      node768 = node767_l;
      node769 = node767_r;
      node770 = node766_r;
      node771 = node765_r;
      node772 = node764_r;
      node773_r = node731_r & pixel[358];
      node773_l = node731_r & ~pixel[358];
      node774_r = node773_l & pixel[267];
      node774_l = node773_l & ~pixel[267];
      node775_r = node774_l & pixel[155];
      node775_l = node774_l & ~pixel[155];
      node776_r = node775_l & pixel[330];
      node776_l = node775_l & ~pixel[330];
      node777_r = node776_l & pixel[378];
      node777_l = node776_l & ~pixel[378];
      node778 = node777_l;
      node779 = node777_r;
      node780 = node776_r;
      node781_r = node775_r & pixel[656];
      node781_l = node775_r & ~pixel[656];
      node782_r = node781_l & pixel[344];
      node782_l = node781_l & ~pixel[344];
      node783 = node782_l;
      node784 = node782_r;
      node785_r = node781_r & pixel[686];
      node785_l = node781_r & ~pixel[686];
      node786 = node785_l;
      node787 = node785_r;
      node788_r = node774_r & pixel[156];
      node788_l = node774_r & ~pixel[156];
      node789_r = node788_l & pixel[631];
      node789_l = node788_l & ~pixel[631];
      node790_r = node789_l & pixel[385];
      node790_l = node789_l & ~pixel[385];
      node791 = node790_l;
      node792 = node790_r;
      node793_r = node789_r & pixel[741];
      node793_l = node789_r & ~pixel[741];
      node794 = node793_l;
      node795 = node793_r;
      node796_r = node788_r & pixel[498];
      node796_l = node788_r & ~pixel[498];
      node797_r = node796_l & pixel[375];
      node797_l = node796_l & ~pixel[375];
      node798 = node797_l;
      node799 = node797_r;
      node800_r = node796_r & pixel[623];
      node800_l = node796_r & ~pixel[623];
      node801 = node800_l;
      node802 = node800_r;
      node803_r = node773_r & pixel[216];
      node803_l = node773_r & ~pixel[216];
      node804_r = node803_l & pixel[243];
      node804_l = node803_l & ~pixel[243];
      node805_r = node804_l & pixel[574];
      node805_l = node804_l & ~pixel[574];
      node806_r = node805_l & pixel[718];
      node806_l = node805_l & ~pixel[718];
      node807 = node806_l;
      node808 = node806_r;
      node809_r = node805_r & pixel[382];
      node809_l = node805_r & ~pixel[382];
      node810 = node809_l;
      node811 = node809_r;
      node812_r = node804_r & pixel[303];
      node812_l = node804_r & ~pixel[303];
      node813_r = node812_l & pixel[681];
      node813_l = node812_l & ~pixel[681];
      node814 = node813_l;
      node815 = node813_r;
      node816_r = node812_r & pixel[242];
      node816_l = node812_r & ~pixel[242];
      node817 = node816_l;
      node818 = node816_r;
      node819_r = node803_r & pixel[626];
      node819_l = node803_r & ~pixel[626];
      node820_r = node819_l & pixel[208];
      node820_l = node819_l & ~pixel[208];
      node821_r = node820_l & pixel[486];
      node821_l = node820_l & ~pixel[486];
      node822 = node821_l;
      node823 = node821_r;
      node824_r = node820_r & pixel[509];
      node824_l = node820_r & ~pixel[509];
      node825 = node824_l;
      node826 = node824_r;
      node827_r = node819_r & pixel[344];
      node827_l = node819_r & ~pixel[344];
      node828_r = node827_l & pixel[708];
      node828_l = node827_l & ~pixel[708];
      node829 = node828_l;
      node830 = node828_r;
      node831_r = node827_r & pixel[710];
      node831_l = node827_r & ~pixel[710];
      node832 = node831_l;
      node833 = node831_r;
      node834_r = node0_r & pixel[263];
      node834_l = node0_r & ~pixel[263];
      node835_r = node834_l & pixel[204];
      node835_l = node834_l & ~pixel[204];
      node836_r = node835_l & pixel[410];
      node836_l = node835_l & ~pixel[410];
      node837_r = node836_l & pixel[577];
      node837_l = node836_l & ~pixel[577];
      node838_r = node837_l & pixel[465];
      node838_l = node837_l & ~pixel[465];
      node839_r = node838_l & pixel[300];
      node839_l = node838_l & ~pixel[300];
      node840_r = node839_l & pixel[374];
      node840_l = node839_l & ~pixel[374];
      node841_r = node840_l & pixel[206];
      node841_l = node840_l & ~pixel[206];
      node842_r = node841_l & pixel[319];
      node842_l = node841_l & ~pixel[319];
      node843 = node842_l;
      node844 = node842_r;
      node845_r = node841_r & pixel[542];
      node845_l = node841_r & ~pixel[542];
      node846 = node845_l;
      node847 = node845_r;
      node848_r = node840_r & pixel[595];
      node848_l = node840_r & ~pixel[595];
      node849_r = node848_l & pixel[352];
      node849_l = node848_l & ~pixel[352];
      node850 = node849_l;
      node851 = node849_r;
      node852_r = node848_r & pixel[132];
      node852_l = node848_r & ~pixel[132];
      node853 = node852_l;
      node854 = node852_r;
      node855_r = node839_r & pixel[654];
      node855_l = node839_r & ~pixel[654];
      node856_r = node855_l & pixel[650];
      node856_l = node855_l & ~pixel[650];
      node857_r = node856_l & pixel[353];
      node857_l = node856_l & ~pixel[353];
      node858 = node857_l;
      node859 = node857_r;
      node860_r = node856_r & pixel[575];
      node860_l = node856_r & ~pixel[575];
      node861 = node860_l;
      node862 = node860_r;
      node863_r = node855_r & pixel[184];
      node863_l = node855_r & ~pixel[184];
      node864_r = node863_l & pixel[239];
      node864_l = node863_l & ~pixel[239];
      node865 = node864_l;
      node866 = node864_r;
      node867_r = node863_r & pixel[265];
      node867_l = node863_r & ~pixel[265];
      node868 = node867_l;
      node869 = node867_r;
      node870_r = node838_r & pixel[248];
      node870_l = node838_r & ~pixel[248];
      node871_r = node870_l & pixel[401];
      node871_l = node870_l & ~pixel[401];
      node872_r = node871_l & pixel[266];
      node872_l = node871_l & ~pixel[266];
      node873_r = node872_l & pixel[496];
      node873_l = node872_l & ~pixel[496];
      node874 = node873_l;
      node875 = node873_r;
      node876_r = node872_r & pixel[654];
      node876_l = node872_r & ~pixel[654];
      node877 = node876_l;
      node878 = node876_r;
      node879_r = node871_r & pixel[484];
      node879_l = node871_r & ~pixel[484];
      node880_r = node879_l & pixel[567];
      node880_l = node879_l & ~pixel[567];
      node881 = node880_l;
      node882 = node880_r;
      node883_r = node879_r & pixel[321];
      node883_l = node879_r & ~pixel[321];
      node884 = node883_l;
      node885 = node883_r;
      node886_r = node870_r & pixel[459];
      node886_l = node870_r & ~pixel[459];
      node887_r = node886_l & pixel[440];
      node887_l = node886_l & ~pixel[440];
      node888 = node887_l;
      node889 = node887_r;
      node890_r = node886_r & pixel[164];
      node890_l = node886_r & ~pixel[164];
      node891_r = node890_l & pixel[492];
      node891_l = node890_l & ~pixel[492];
      node892 = node891_l;
      node893 = node891_r;
      node894 = node890_r;
      node895_r = node837_r & pixel[656];
      node895_l = node837_r & ~pixel[656];
      node896_r = node895_l & pixel[660];
      node896_l = node895_l & ~pixel[660];
      node897_r = node896_l & pixel[513];
      node897_l = node896_l & ~pixel[513];
      node898_r = node897_l & pixel[347];
      node898_l = node897_l & ~pixel[347];
      node899_r = node898_l & pixel[516];
      node899_l = node898_l & ~pixel[516];
      node900 = node899_l;
      node901 = node899_r;
      node902_r = node898_r & pixel[346];
      node902_l = node898_r & ~pixel[346];
      node903 = node902_l;
      node904 = node902_r;
      node905_r = node897_r & pixel[465];
      node905_l = node897_r & ~pixel[465];
      node906_r = node905_l & pixel[319];
      node906_l = node905_l & ~pixel[319];
      node907 = node906_l;
      node908 = node906_r;
      node909_r = node905_r & pixel[607];
      node909_l = node905_r & ~pixel[607];
      node910 = node909_l;
      node911 = node909_r;
      node912_r = node896_r & pixel[353];
      node912_l = node896_r & ~pixel[353];
      node913_r = node912_l & pixel[579];
      node913_l = node912_l & ~pixel[579];
      node914_r = node913_l & pixel[346];
      node914_l = node913_l & ~pixel[346];
      node915 = node914_l;
      node916 = node914_r;
      node917_r = node913_r & pixel[519];
      node917_l = node913_r & ~pixel[519];
      node918 = node917_l;
      node919 = node917_r;
      node920_r = node912_r & pixel[508];
      node920_l = node912_r & ~pixel[508];
      node921_r = node920_l & pixel[711];
      node921_l = node920_l & ~pixel[711];
      node922 = node921_l;
      node923 = node921_r;
      node924 = node920_r;
      node925_r = node895_r & pixel[262];
      node925_l = node895_r & ~pixel[262];
      node926_r = node925_l & pixel[293];
      node926_l = node925_l & ~pixel[293];
      node927_r = node926_l & pixel[492];
      node927_l = node926_l & ~pixel[492];
      node928_r = node927_l & pixel[523];
      node928_l = node927_l & ~pixel[523];
      node929 = node928_l;
      node930 = node928_r;
      node931_r = node927_r & pixel[317];
      node931_l = node927_r & ~pixel[317];
      node932 = node931_l;
      node933 = node931_r;
      node934_r = node926_r & pixel[205];
      node934_l = node926_r & ~pixel[205];
      node935_r = node934_l & pixel[178];
      node935_l = node934_l & ~pixel[178];
      node936 = node935_l;
      node937 = node935_r;
      node938 = node934_r;
      node939_r = node925_r & pixel[483];
      node939_l = node925_r & ~pixel[483];
      node940_r = node939_l & pixel[380];
      node940_l = node939_l & ~pixel[380];
      node941_r = node940_l & pixel[716];
      node941_l = node940_l & ~pixel[716];
      node942 = node941_l;
      node943 = node941_r;
      node944_r = node940_r & pixel[347];
      node944_l = node940_r & ~pixel[347];
      node945 = node944_l;
      node946 = node944_r;
      node947_r = node939_r & pixel[601];
      node947_l = node939_r & ~pixel[601];
      node948 = node947_l;
      node949_r = node947_r & pixel[327];
      node949_l = node947_r & ~pixel[327];
      node950 = node949_l;
      node951 = node949_r;
      node952_r = node836_r & pixel[153];
      node952_l = node836_r & ~pixel[153];
      node953_r = node952_l & pixel[266];
      node953_l = node952_l & ~pixel[266];
      node954_r = node953_l & pixel[514];
      node954_l = node953_l & ~pixel[514];
      node955_r = node954_l & pixel[595];
      node955_l = node954_l & ~pixel[595];
      node956_r = node955_l & pixel[210];
      node956_l = node955_l & ~pixel[210];
      node957_r = node956_l & pixel[538];
      node957_l = node956_l & ~pixel[538];
      node958 = node957_l;
      node959 = node957_r;
      node960_r = node956_r & pixel[653];
      node960_l = node956_r & ~pixel[653];
      node961 = node960_l;
      node962 = node960_r;
      node963_r = node955_r & pixel[377];
      node963_l = node955_r & ~pixel[377];
      node964 = node963_l;
      node965_r = node963_r & pixel[483];
      node965_l = node963_r & ~pixel[483];
      node966 = node965_l;
      node967 = node965_r;
      node968_r = node954_r & pixel[625];
      node968_l = node954_r & ~pixel[625];
      node969_r = node968_l & pixel[483];
      node969_l = node968_l & ~pixel[483];
      node970_r = node969_l & pixel[122];
      node970_l = node969_l & ~pixel[122];
      node971 = node970_l;
      node972 = node970_r;
      node973_r = node969_r & pixel[415];
      node973_l = node969_r & ~pixel[415];
      node974 = node973_l;
      node975 = node973_r;
      node976_r = node968_r & pixel[536];
      node976_l = node968_r & ~pixel[536];
      node977_r = node976_l & pixel[181];
      node977_l = node976_l & ~pixel[181];
      node978 = node977_l;
      node979 = node977_r;
      node980_r = node976_r & pixel[547];
      node980_l = node976_r & ~pixel[547];
      node981 = node980_l;
      node982 = node980_r;
      node983_r = node953_r & pixel[242];
      node983_l = node953_r & ~pixel[242];
      node984_r = node983_l & pixel[655];
      node984_l = node983_l & ~pixel[655];
      node985_r = node984_l & pixel[574];
      node985_l = node984_l & ~pixel[574];
      node986_r = node985_l & pixel[514];
      node986_l = node985_l & ~pixel[514];
      node987 = node986_l;
      node988 = node986_r;
      node989_r = node985_r & pixel[273];
      node989_l = node985_r & ~pixel[273];
      node990 = node989_l;
      node991 = node989_r;
      node992_r = node984_r & pixel[566];
      node992_l = node984_r & ~pixel[566];
      node993_r = node992_l & pixel[483];
      node993_l = node992_l & ~pixel[483];
      node994 = node993_l;
      node995 = node993_r;
      node996_r = node992_r & pixel[493];
      node996_l = node992_r & ~pixel[493];
      node997 = node996_l;
      node998 = node996_r;
      node999_r = node983_r & pixel[325];
      node999_l = node983_r & ~pixel[325];
      node1000_r = node999_l & pixel[245];
      node1000_l = node999_l & ~pixel[245];
      node1001_r = node1000_l & pixel[296];
      node1001_l = node1000_l & ~pixel[296];
      node1002 = node1001_l;
      node1003 = node1001_r;
      node1004_r = node1000_r & pixel[328];
      node1004_l = node1000_r & ~pixel[328];
      node1005 = node1004_l;
      node1006 = node1004_r;
      node1007_r = node999_r & pixel[511];
      node1007_l = node999_r & ~pixel[511];
      node1008_r = node1007_l & pixel[411];
      node1008_l = node1007_l & ~pixel[411];
      node1009 = node1008_l;
      node1010 = node1008_r;
      node1011_r = node1007_r & pixel[209];
      node1011_l = node1007_r & ~pixel[209];
      node1012 = node1011_l;
      node1013 = node1011_r;
      node1014_r = node952_r & pixel[296];
      node1014_l = node952_r & ~pixel[296];
      node1015_r = node1014_l & pixel[658];
      node1015_l = node1014_l & ~pixel[658];
      node1016_r = node1015_l & pixel[540];
      node1016_l = node1015_l & ~pixel[540];
      node1017_r = node1016_l & pixel[567];
      node1017_l = node1016_l & ~pixel[567];
      node1018_r = node1017_l & pixel[626];
      node1018_l = node1017_l & ~pixel[626];
      node1019 = node1018_l;
      node1020 = node1018_r;
      node1021_r = node1017_r & pixel[352];
      node1021_l = node1017_r & ~pixel[352];
      node1022 = node1021_l;
      node1023 = node1021_r;
      node1024_r = node1016_r & pixel[290];
      node1024_l = node1016_r & ~pixel[290];
      node1025_r = node1024_l & pixel[429];
      node1025_l = node1024_l & ~pixel[429];
      node1026 = node1025_l;
      node1027 = node1025_r;
      node1028_r = node1024_r & pixel[456];
      node1028_l = node1024_r & ~pixel[456];
      node1029 = node1028_l;
      node1030 = node1028_r;
      node1031_r = node1015_r & pixel[290];
      node1031_l = node1015_r & ~pixel[290];
      node1032_r = node1031_l & pixel[123];
      node1032_l = node1031_l & ~pixel[123];
      node1033_r = node1032_l & pixel[661];
      node1033_l = node1032_l & ~pixel[661];
      node1034 = node1033_l;
      node1035 = node1033_r;
      node1036_r = node1032_r & pixel[485];
      node1036_l = node1032_r & ~pixel[485];
      node1037 = node1036_l;
      node1038 = node1036_r;
      node1039_r = node1031_r & pixel[326];
      node1039_l = node1031_r & ~pixel[326];
      node1040_r = node1039_l & pixel[487];
      node1040_l = node1039_l & ~pixel[487];
      node1041 = node1040_l;
      node1042 = node1040_r;
      node1043_r = node1039_r & pixel[434];
      node1043_l = node1039_r & ~pixel[434];
      node1044 = node1043_l;
      node1045 = node1043_r;
      node1046_r = node1014_r & pixel[488];
      node1046_l = node1014_r & ~pixel[488];
      node1047_r = node1046_l & pixel[513];
      node1047_l = node1046_l & ~pixel[513];
      node1048_r = node1047_l & pixel[91];
      node1048_l = node1047_l & ~pixel[91];
      node1049_r = node1048_l & pixel[348];
      node1049_l = node1048_l & ~pixel[348];
      node1050 = node1049_l;
      node1051 = node1049_r;
      node1052_r = node1048_r & pixel[612];
      node1052_l = node1048_r & ~pixel[612];
      node1053 = node1052_l;
      node1054 = node1052_r;
      node1055_r = node1047_r & pixel[456];
      node1055_l = node1047_r & ~pixel[456];
      node1056_r = node1055_l & pixel[600];
      node1056_l = node1055_l & ~pixel[600];
      node1057 = node1056_l;
      node1058 = node1056_r;
      node1059_r = node1055_r & pixel[594];
      node1059_l = node1055_r & ~pixel[594];
      node1060 = node1059_l;
      node1061 = node1059_r;
      node1062_r = node1046_r & pixel[233];
      node1062_l = node1046_r & ~pixel[233];
      node1063_r = node1062_l & pixel[322];
      node1063_l = node1062_l & ~pixel[322];
      node1064_r = node1063_l & pixel[685];
      node1064_l = node1063_l & ~pixel[685];
      node1065 = node1064_l;
      node1066 = node1064_r;
      node1067_r = node1063_r & pixel[550];
      node1067_l = node1063_r & ~pixel[550];
      node1068 = node1067_l;
      node1069 = node1067_r;
      node1070_r = node1062_r & pixel[289];
      node1070_l = node1062_r & ~pixel[289];
      node1071_r = node1070_l & pixel[489];
      node1071_l = node1070_l & ~pixel[489];
      node1072 = node1071_l;
      node1073 = node1071_r;
      node1074_r = node1070_r & pixel[664];
      node1074_l = node1070_r & ~pixel[664];
      node1075 = node1074_l;
      node1076 = node1074_r;
      node1077_r = node835_r & pixel[517];
      node1077_l = node835_r & ~pixel[517];
      node1078_r = node1077_l & pixel[370];
      node1078_l = node1077_l & ~pixel[370];
      node1079_r = node1078_l & pixel[290];
      node1079_l = node1078_l & ~pixel[290];
      node1080_r = node1079_l & pixel[546];
      node1080_l = node1079_l & ~pixel[546];
      node1081_r = node1080_l & pixel[513];
      node1081_l = node1080_l & ~pixel[513];
      node1082_r = node1081_l & pixel[180];
      node1082_l = node1081_l & ~pixel[180];
      node1083_r = node1082_l & pixel[321];
      node1083_l = node1082_l & ~pixel[321];
      node1084 = node1083_l;
      node1085 = node1083_r;
      node1086_r = node1082_r & pixel[515];
      node1086_l = node1082_r & ~pixel[515];
      node1087 = node1086_l;
      node1088 = node1086_r;
      node1089_r = node1081_r & pixel[486];
      node1089_l = node1081_r & ~pixel[486];
      node1090_r = node1089_l & pixel[343];
      node1090_l = node1089_l & ~pixel[343];
      node1091 = node1090_l;
      node1092 = node1090_r;
      node1093_r = node1089_r & pixel[373];
      node1093_l = node1089_r & ~pixel[373];
      node1094 = node1093_l;
      node1095 = node1093_r;
      node1096_r = node1080_r & pixel[514];
      node1096_l = node1080_r & ~pixel[514];
      node1097_r = node1096_l & pixel[209];
      node1097_l = node1096_l & ~pixel[209];
      node1098_r = node1097_l & pixel[154];
      node1098_l = node1097_l & ~pixel[154];
      node1099 = node1098_l;
      node1100 = node1098_r;
      node1101_r = node1097_r & pixel[455];
      node1101_l = node1097_r & ~pixel[455];
      node1102 = node1101_l;
      node1103 = node1101_r;
      node1104_r = node1096_r & pixel[228];
      node1104_l = node1096_r & ~pixel[228];
      node1105_r = node1104_l & pixel[374];
      node1105_l = node1104_l & ~pixel[374];
      node1106 = node1105_l;
      node1107 = node1105_r;
      node1108 = node1104_r;
      node1109_r = node1079_r & pixel[183];
      node1109_l = node1079_r & ~pixel[183];
      node1110_r = node1109_l & pixel[570];
      node1110_l = node1109_l & ~pixel[570];
      node1111_r = node1110_l & pixel[181];
      node1111_l = node1110_l & ~pixel[181];
      node1112_r = node1111_l & pixel[66];
      node1112_l = node1111_l & ~pixel[66];
      node1113 = node1112_l;
      node1114 = node1112_r;
      node1115_r = node1111_r & pixel[151];
      node1115_l = node1111_r & ~pixel[151];
      node1116 = node1115_l;
      node1117 = node1115_r;
      node1118_r = node1110_r & pixel[628];
      node1118_l = node1110_r & ~pixel[628];
      node1119_r = node1118_l & pixel[526];
      node1119_l = node1118_l & ~pixel[526];
      node1120 = node1119_l;
      node1121 = node1119_r;
      node1122_r = node1118_r & pixel[595];
      node1122_l = node1118_r & ~pixel[595];
      node1123 = node1122_l;
      node1124 = node1122_r;
      node1125_r = node1109_r & pixel[514];
      node1125_l = node1109_r & ~pixel[514];
      node1126_r = node1125_l & pixel[267];
      node1126_l = node1125_l & ~pixel[267];
      node1127_r = node1126_l & pixel[234];
      node1127_l = node1126_l & ~pixel[234];
      node1128 = node1127_l;
      node1129 = node1127_r;
      node1130_r = node1126_r & pixel[209];
      node1130_l = node1126_r & ~pixel[209];
      node1131 = node1130_l;
      node1132 = node1130_r;
      node1133_r = node1125_r & pixel[612];
      node1133_l = node1125_r & ~pixel[612];
      node1134_r = node1133_l & pixel[289];
      node1134_l = node1133_l & ~pixel[289];
      node1135 = node1134_l;
      node1136 = node1134_r;
      node1137 = node1133_r;
      node1138_r = node1078_r & pixel[181];
      node1138_l = node1078_r & ~pixel[181];
      node1139_r = node1138_l & pixel[121];
      node1139_l = node1138_l & ~pixel[121];
      node1140_r = node1139_l & pixel[90];
      node1140_l = node1139_l & ~pixel[90];
      node1141_r = node1140_l & pixel[437];
      node1141_l = node1140_l & ~pixel[437];
      node1142_r = node1141_l & pixel[542];
      node1142_l = node1141_l & ~pixel[542];
      node1143 = node1142_l;
      node1144 = node1142_r;
      node1145_r = node1141_r & pixel[237];
      node1145_l = node1141_r & ~pixel[237];
      node1146 = node1145_l;
      node1147 = node1145_r;
      node1148 = node1140_r;
      node1149_r = node1139_r & pixel[431];
      node1149_l = node1139_r & ~pixel[431];
      node1150_r = node1149_l & pixel[157];
      node1150_l = node1149_l & ~pixel[157];
      node1151 = node1150_l;
      node1152 = node1150_r;
      node1153_r = node1149_r & pixel[124];
      node1153_l = node1149_r & ~pixel[124];
      node1154_r = node1153_l & pixel[355];
      node1154_l = node1153_l & ~pixel[355];
      node1155 = node1154_l;
      node1156 = node1154_r;
      node1157_r = node1153_r & pixel[528];
      node1157_l = node1153_r & ~pixel[528];
      node1158 = node1157_l;
      node1159 = node1157_r;
      node1160_r = node1138_r & pixel[526];
      node1160_l = node1138_r & ~pixel[526];
      node1161_r = node1160_l & pixel[629];
      node1161_l = node1160_l & ~pixel[629];
      node1162_r = node1161_l & pixel[653];
      node1162_l = node1161_l & ~pixel[653];
      node1163_r = node1162_l & pixel[683];
      node1163_l = node1162_l & ~pixel[683];
      node1164 = node1163_l;
      node1165 = node1163_r;
      node1166_r = node1162_r & pixel[630];
      node1166_l = node1162_r & ~pixel[630];
      node1167 = node1166_l;
      node1168 = node1166_r;
      node1169_r = node1161_r & pixel[301];
      node1169_l = node1161_r & ~pixel[301];
      node1170_r = node1169_l & pixel[466];
      node1170_l = node1169_l & ~pixel[466];
      node1171 = node1170_l;
      node1172 = node1170_r;
      node1173_r = node1169_r & pixel[607];
      node1173_l = node1169_r & ~pixel[607];
      node1174 = node1173_l;
      node1175 = node1173_r;
      node1176_r = node1160_r & pixel[322];
      node1176_l = node1160_r & ~pixel[322];
      node1177_r = node1176_l & pixel[98];
      node1177_l = node1176_l & ~pixel[98];
      node1178_r = node1177_l & pixel[512];
      node1178_l = node1177_l & ~pixel[512];
      node1179 = node1178_l;
      node1180 = node1178_r;
      node1181 = node1177_r;
      node1182_r = node1176_r & pixel[512];
      node1182_l = node1176_r & ~pixel[512];
      node1183_r = node1182_l & pixel[658];
      node1183_l = node1182_l & ~pixel[658];
      node1184 = node1183_l;
      node1185 = node1183_r;
      node1186_r = node1182_r & pixel[175];
      node1186_l = node1182_r & ~pixel[175];
      node1187 = node1186_l;
      node1188 = node1186_r;
      node1189_r = node1077_r & pixel[400];
      node1189_l = node1077_r & ~pixel[400];
      node1190_r = node1189_l & pixel[582];
      node1190_l = node1189_l & ~pixel[582];
      node1191_r = node1190_l & pixel[660];
      node1191_l = node1190_l & ~pixel[660];
      node1192_r = node1191_l & pixel[597];
      node1192_l = node1191_l & ~pixel[597];
      node1193_r = node1192_l & pixel[542];
      node1193_l = node1192_l & ~pixel[542];
      node1194_r = node1193_l & pixel[149];
      node1194_l = node1193_l & ~pixel[149];
      node1195 = node1194_l;
      node1196 = node1194_r;
      node1197_r = node1193_r & pixel[359];
      node1197_l = node1193_r & ~pixel[359];
      node1198 = node1197_l;
      node1199 = node1197_r;
      node1200_r = node1192_r & pixel[345];
      node1200_l = node1192_r & ~pixel[345];
      node1201_r = node1200_l & pixel[426];
      node1201_l = node1200_l & ~pixel[426];
      node1202 = node1201_l;
      node1203 = node1201_r;
      node1204_r = node1200_r & pixel[462];
      node1204_l = node1200_r & ~pixel[462];
      node1205 = node1204_l;
      node1206 = node1204_r;
      node1207_r = node1191_r & pixel[346];
      node1207_l = node1191_r & ~pixel[346];
      node1208_r = node1207_l & pixel[154];
      node1208_l = node1207_l & ~pixel[154];
      node1209_r = node1208_l & pixel[574];
      node1209_l = node1208_l & ~pixel[574];
      node1210 = node1209_l;
      node1211 = node1209_r;
      node1212_r = node1208_r & pixel[549];
      node1212_l = node1208_r & ~pixel[549];
      node1213 = node1212_l;
      node1214 = node1212_r;
      node1215_r = node1207_r & pixel[432];
      node1215_l = node1207_r & ~pixel[432];
      node1216_r = node1215_l & pixel[634];
      node1216_l = node1215_l & ~pixel[634];
      node1217 = node1216_l;
      node1218 = node1216_r;
      node1219_r = node1215_r & pixel[629];
      node1219_l = node1215_r & ~pixel[629];
      node1220 = node1219_l;
      node1221 = node1219_r;
      node1222_r = node1190_r & pixel[386];
      node1222_l = node1190_r & ~pixel[386];
      node1223_r = node1222_l & pixel[690];
      node1223_l = node1222_l & ~pixel[690];
      node1224_r = node1223_l & pixel[375];
      node1224_l = node1223_l & ~pixel[375];
      node1225_r = node1224_l & pixel[657];
      node1225_l = node1224_l & ~pixel[657];
      node1226 = node1225_l;
      node1227 = node1225_r;
      node1228_r = node1224_r & pixel[550];
      node1228_l = node1224_r & ~pixel[550];
      node1229 = node1228_l;
      node1230 = node1228_r;
      node1231_r = node1223_r & pixel[348];
      node1231_l = node1223_r & ~pixel[348];
      node1232 = node1231_l;
      node1233 = node1231_r;
      node1234_r = node1222_r & pixel[369];
      node1234_l = node1222_r & ~pixel[369];
      node1235_r = node1234_l & pixel[382];
      node1235_l = node1234_l & ~pixel[382];
      node1236 = node1235_l;
      node1237_r = node1235_r & pixel[185];
      node1237_l = node1235_r & ~pixel[185];
      node1238 = node1237_l;
      node1239 = node1237_r;
      node1240 = node1234_r;
      node1241_r = node1189_r & pixel[657];
      node1241_l = node1189_r & ~pixel[657];
      node1242_r = node1241_l & pixel[182];
      node1242_l = node1241_l & ~pixel[182];
      node1243_r = node1242_l & pixel[150];
      node1243_l = node1242_l & ~pixel[150];
      node1244_r = node1243_l & pixel[382];
      node1244_l = node1243_l & ~pixel[382];
      node1245_r = node1244_l & pixel[575];
      node1245_l = node1244_l & ~pixel[575];
      node1246 = node1245_l;
      node1247 = node1245_r;
      node1248_r = node1244_r & pixel[498];
      node1248_l = node1244_r & ~pixel[498];
      node1249 = node1248_l;
      node1250 = node1248_r;
      node1251_r = node1243_r & pixel[316];
      node1251_l = node1243_r & ~pixel[316];
      node1252_r = node1251_l & pixel[370];
      node1252_l = node1251_l & ~pixel[370];
      node1253 = node1252_l;
      node1254 = node1252_r;
      node1255_r = node1251_r & pixel[239];
      node1255_l = node1251_r & ~pixel[239];
      node1256 = node1255_l;
      node1257 = node1255_r;
      node1258_r = node1242_r & pixel[287];
      node1258_l = node1242_r & ~pixel[287];
      node1259_r = node1258_l & pixel[687];
      node1259_l = node1258_l & ~pixel[687];
      node1260_r = node1259_l & pixel[681];
      node1260_l = node1259_l & ~pixel[681];
      node1261 = node1260_l;
      node1262 = node1260_r;
      node1263 = node1259_r;
      node1264_r = node1258_r & pixel[661];
      node1264_l = node1258_r & ~pixel[661];
      node1265_r = node1264_l & pixel[543];
      node1265_l = node1264_l & ~pixel[543];
      node1266 = node1265_l;
      node1267 = node1265_r;
      node1268_r = node1264_r & pixel[241];
      node1268_l = node1264_r & ~pixel[241];
      node1269 = node1268_l;
      node1270 = node1268_r;
      node1271_r = node1241_r & pixel[183];
      node1271_l = node1241_r & ~pixel[183];
      node1272_r = node1271_l & pixel[381];
      node1272_l = node1271_l & ~pixel[381];
      node1273 = node1272_l;
      node1274 = node1272_r;
      node1275_r = node1271_r & pixel[371];
      node1275_l = node1271_r & ~pixel[371];
      node1276_r = node1275_l & pixel[432];
      node1276_l = node1275_l & ~pixel[432];
      node1277 = node1276_l;
      node1278_r = node1276_r & pixel[485];
      node1278_l = node1276_r & ~pixel[485];
      node1279 = node1278_l;
      node1280 = node1278_r;
      node1281_r = node1275_r & pixel[173];
      node1281_l = node1275_r & ~pixel[173];
      node1282_r = node1281_l & pixel[470];
      node1282_l = node1281_l & ~pixel[470];
      node1283 = node1282_l;
      node1284 = node1282_r;
      node1285_r = node1281_r & pixel[442];
      node1285_l = node1281_r & ~pixel[442];
      node1286 = node1285_l;
      node1287 = node1285_r;
      node1288_r = node834_r & pixel[158];
      node1288_l = node834_r & ~pixel[158];
      node1289_r = node1288_l & pixel[98];
      node1289_l = node1288_l & ~pixel[98];
      node1290_r = node1289_l & pixel[713];
      node1290_l = node1289_l & ~pixel[713];
      node1291_r = node1290_l & pixel[239];
      node1291_l = node1290_l & ~pixel[239];
      node1292_r = node1291_l & pixel[153];
      node1292_l = node1291_l & ~pixel[153];
      node1293_r = node1292_l & pixel[211];
      node1293_l = node1292_l & ~pixel[211];
      node1294_r = node1293_l & pixel[67];
      node1294_l = node1293_l & ~pixel[67];
      node1295_r = node1294_l & pixel[327];
      node1295_l = node1294_l & ~pixel[327];
      node1296 = node1295_l;
      node1297 = node1295_r;
      node1298 = node1294_r;
      node1299_r = node1293_r & pixel[571];
      node1299_l = node1293_r & ~pixel[571];
      node1300_r = node1299_l & pixel[349];
      node1300_l = node1299_l & ~pixel[349];
      node1301 = node1300_l;
      node1302 = node1300_r;
      node1303_r = node1299_r & pixel[495];
      node1303_l = node1299_r & ~pixel[495];
      node1304 = node1303_l;
      node1305 = node1303_r;
      node1306_r = node1292_r & pixel[628];
      node1306_l = node1292_r & ~pixel[628];
      node1307_r = node1306_l & pixel[322];
      node1307_l = node1306_l & ~pixel[322];
      node1308_r = node1307_l & pixel[97];
      node1308_l = node1307_l & ~pixel[97];
      node1309 = node1308_l;
      node1310 = node1308_r;
      node1311_r = node1307_r & pixel[459];
      node1311_l = node1307_r & ~pixel[459];
      node1312 = node1311_l;
      node1313 = node1311_r;
      node1314_r = node1306_r & pixel[399];
      node1314_l = node1306_r & ~pixel[399];
      node1315_r = node1314_l & pixel[374];
      node1315_l = node1314_l & ~pixel[374];
      node1316 = node1315_l;
      node1317 = node1315_r;
      node1318_r = node1314_r & pixel[605];
      node1318_l = node1314_r & ~pixel[605];
      node1319 = node1318_l;
      node1320 = node1318_r;
      node1321_r = node1291_r & pixel[381];
      node1321_l = node1291_r & ~pixel[381];
      node1322_r = node1321_l & pixel[272];
      node1322_l = node1321_l & ~pixel[272];
      node1323_r = node1322_l & pixel[189];
      node1323_l = node1322_l & ~pixel[189];
      node1324_r = node1323_l & pixel[544];
      node1324_l = node1323_l & ~pixel[544];
      node1325 = node1324_l;
      node1326 = node1324_r;
      node1327_r = node1323_r & pixel[516];
      node1327_l = node1323_r & ~pixel[516];
      node1328 = node1327_l;
      node1329 = node1327_r;
      node1330_r = node1322_r & pixel[344];
      node1330_l = node1322_r & ~pixel[344];
      node1331_r = node1330_l & pixel[326];
      node1331_l = node1330_l & ~pixel[326];
      node1332 = node1331_l;
      node1333 = node1331_r;
      node1334_r = node1330_r & pixel[388];
      node1334_l = node1330_r & ~pixel[388];
      node1335 = node1334_l;
      node1336 = node1334_r;
      node1337_r = node1321_r & pixel[718];
      node1337_l = node1321_r & ~pixel[718];
      node1338_r = node1337_l & pixel[152];
      node1338_l = node1337_l & ~pixel[152];
      node1339_r = node1338_l & pixel[542];
      node1339_l = node1338_l & ~pixel[542];
      node1340 = node1339_l;
      node1341 = node1339_r;
      node1342_r = node1338_r & pixel[515];
      node1342_l = node1338_r & ~pixel[515];
      node1343 = node1342_l;
      node1344 = node1342_r;
      node1345_r = node1337_r & pixel[574];
      node1345_l = node1337_r & ~pixel[574];
      node1346_r = node1345_l & pixel[443];
      node1346_l = node1345_l & ~pixel[443];
      node1347 = node1346_l;
      node1348 = node1346_r;
      node1349_r = node1345_r & pixel[203];
      node1349_l = node1345_r & ~pixel[203];
      node1350 = node1349_l;
      node1351 = node1349_r;
      node1352_r = node1290_r & pixel[317];
      node1352_l = node1290_r & ~pixel[317];
      node1353_r = node1352_l & pixel[204];
      node1353_l = node1352_l & ~pixel[204];
      node1354_r = node1353_l & pixel[601];
      node1354_l = node1353_l & ~pixel[601];
      node1355_r = node1354_l & pixel[600];
      node1355_l = node1354_l & ~pixel[600];
      node1356_r = node1355_l & pixel[266];
      node1356_l = node1355_l & ~pixel[266];
      node1357 = node1356_l;
      node1358 = node1356_r;
      node1359_r = node1355_r & pixel[569];
      node1359_l = node1355_r & ~pixel[569];
      node1360 = node1359_l;
      node1361 = node1359_r;
      node1362_r = node1354_r & pixel[377];
      node1362_l = node1354_r & ~pixel[377];
      node1363_r = node1362_l & pixel[373];
      node1363_l = node1362_l & ~pixel[373];
      node1364 = node1363_l;
      node1365 = node1363_r;
      node1366_r = node1362_r & pixel[433];
      node1366_l = node1362_r & ~pixel[433];
      node1367 = node1366_l;
      node1368 = node1366_r;
      node1369_r = node1353_r & pixel[489];
      node1369_l = node1353_r & ~pixel[489];
      node1370_r = node1369_l & pixel[181];
      node1370_l = node1369_l & ~pixel[181];
      node1371_r = node1370_l & pixel[634];
      node1371_l = node1370_l & ~pixel[634];
      node1372 = node1371_l;
      node1373 = node1371_r;
      node1374_r = node1370_r & pixel[350];
      node1374_l = node1370_r & ~pixel[350];
      node1375 = node1374_l;
      node1376 = node1374_r;
      node1377_r = node1369_r & pixel[634];
      node1377_l = node1369_r & ~pixel[634];
      node1378_r = node1377_l & pixel[302];
      node1378_l = node1377_l & ~pixel[302];
      node1379 = node1378_l;
      node1380 = node1378_r;
      node1381_r = node1377_r & pixel[576];
      node1381_l = node1377_r & ~pixel[576];
      node1382 = node1381_l;
      node1383 = node1381_r;
      node1384_r = node1352_r & pixel[212];
      node1384_l = node1352_r & ~pixel[212];
      node1385_r = node1384_l & pixel[740];
      node1385_l = node1384_l & ~pixel[740];
      node1386_r = node1385_l & pixel[238];
      node1386_l = node1385_l & ~pixel[238];
      node1387_r = node1386_l & pixel[295];
      node1387_l = node1386_l & ~pixel[295];
      node1388 = node1387_l;
      node1389 = node1387_r;
      node1390_r = node1386_r & pixel[545];
      node1390_l = node1386_r & ~pixel[545];
      node1391 = node1390_l;
      node1392 = node1390_r;
      node1393_r = node1385_r & pixel[434];
      node1393_l = node1385_r & ~pixel[434];
      node1394 = node1393_l;
      node1395_r = node1393_r & pixel[404];
      node1395_l = node1393_r & ~pixel[404];
      node1396 = node1395_l;
      node1397 = node1395_r;
      node1398_r = node1384_r & pixel[626];
      node1398_l = node1384_r & ~pixel[626];
      node1399_r = node1398_l & pixel[354];
      node1399_l = node1398_l & ~pixel[354];
      node1400_r = node1399_l & pixel[490];
      node1400_l = node1399_l & ~pixel[490];
      node1401 = node1400_l;
      node1402 = node1400_r;
      node1403_r = node1399_r & pixel[571];
      node1403_l = node1399_r & ~pixel[571];
      node1404 = node1403_l;
      node1405 = node1403_r;
      node1406_r = node1398_r & pixel[659];
      node1406_l = node1398_r & ~pixel[659];
      node1407_r = node1406_l & pixel[491];
      node1407_l = node1406_l & ~pixel[491];
      node1408 = node1407_l;
      node1409 = node1407_r;
      node1410_r = node1406_r & pixel[517];
      node1410_l = node1406_r & ~pixel[517];
      node1411 = node1410_l;
      node1412 = node1410_r;
      node1413_r = node1289_r & pixel[626];
      node1413_l = node1289_r & ~pixel[626];
      node1414_r = node1413_l & pixel[242];
      node1414_l = node1413_l & ~pixel[242];
      node1415_r = node1414_l & pixel[268];
      node1415_l = node1414_l & ~pixel[268];
      node1416_r = node1415_l & pixel[487];
      node1416_l = node1415_l & ~pixel[487];
      node1417_r = node1416_l & pixel[548];
      node1417_l = node1416_l & ~pixel[548];
      node1418_r = node1417_l & pixel[400];
      node1418_l = node1417_l & ~pixel[400];
      node1419 = node1418_l;
      node1420 = node1418_r;
      node1421_r = node1417_r & pixel[266];
      node1421_l = node1417_r & ~pixel[266];
      node1422 = node1421_l;
      node1423 = node1421_r;
      node1424_r = node1416_r & pixel[460];
      node1424_l = node1416_r & ~pixel[460];
      node1425_r = node1424_l & pixel[377];
      node1425_l = node1424_l & ~pixel[377];
      node1426 = node1425_l;
      node1427 = node1425_r;
      node1428 = node1424_r;
      node1429_r = node1415_r & pixel[547];
      node1429_l = node1415_r & ~pixel[547];
      node1430_r = node1429_l & pixel[101];
      node1430_l = node1429_l & ~pixel[101];
      node1431 = node1430_l;
      node1432 = node1430_r;
      node1433_r = node1429_r & pixel[212];
      node1433_l = node1429_r & ~pixel[212];
      node1434 = node1433_l;
      node1435_r = node1433_r & pixel[541];
      node1435_l = node1433_r & ~pixel[541];
      node1436 = node1435_l;
      node1437 = node1435_r;
      node1438_r = node1414_r & pixel[345];
      node1438_l = node1414_r & ~pixel[345];
      node1439 = node1438_l;
      node1440 = node1438_r;
      node1441_r = node1413_r & pixel[297];
      node1441_l = node1413_r & ~pixel[297];
      node1442_r = node1441_l & pixel[384];
      node1442_l = node1441_l & ~pixel[384];
      node1443_r = node1442_l & pixel[267];
      node1443_l = node1442_l & ~pixel[267];
      node1444_r = node1443_l & pixel[461];
      node1444_l = node1443_l & ~pixel[461];
      node1445_r = node1444_l & pixel[402];
      node1445_l = node1444_l & ~pixel[402];
      node1446 = node1445_l;
      node1447 = node1445_r;
      node1448 = node1444_r;
      node1449_r = node1443_r & pixel[177];
      node1449_l = node1443_r & ~pixel[177];
      node1450_r = node1449_l & pixel[440];
      node1450_l = node1449_l & ~pixel[440];
      node1451 = node1450_l;
      node1452 = node1450_r;
      node1453 = node1449_r;
      node1454_r = node1442_r & pixel[379];
      node1454_l = node1442_r & ~pixel[379];
      node1455_r = node1454_l & pixel[512];
      node1455_l = node1454_l & ~pixel[512];
      node1456 = node1455_l;
      node1457 = node1455_r;
      node1458 = node1454_r;
      node1459_r = node1441_r & pixel[268];
      node1459_l = node1441_r & ~pixel[268];
      node1460_r = node1459_l & pixel[318];
      node1460_l = node1459_l & ~pixel[318];
      node1461_r = node1460_l & pixel[415];
      node1461_l = node1460_l & ~pixel[415];
      node1462 = node1461_l;
      node1463 = node1461_r;
      node1464 = node1460_r;
      node1465_r = node1459_r & pixel[495];
      node1465_l = node1459_r & ~pixel[495];
      node1466 = node1465_l;
      node1467_r = node1465_r & pixel[357];
      node1467_l = node1465_r & ~pixel[357];
      node1468 = node1467_l;
      node1469 = node1467_r;
      node1470_r = node1288_r & pixel[524];
      node1470_l = node1288_r & ~pixel[524];
      node1471_r = node1470_l & pixel[609];
      node1471_l = node1470_l & ~pixel[609];
      node1472_r = node1471_l & pixel[298];
      node1472_l = node1471_l & ~pixel[298];
      node1473_r = node1472_l & pixel[352];
      node1473_l = node1472_l & ~pixel[352];
      node1474_r = node1473_l & pixel[381];
      node1474_l = node1473_l & ~pixel[381];
      node1475_r = node1474_l & pixel[489];
      node1475_l = node1474_l & ~pixel[489];
      node1476_r = node1475_l & pixel[386];
      node1476_l = node1475_l & ~pixel[386];
      node1477 = node1476_l;
      node1478 = node1476_r;
      node1479_r = node1475_r & pixel[431];
      node1479_l = node1475_r & ~pixel[431];
      node1480 = node1479_l;
      node1481 = node1479_r;
      node1482_r = node1474_r & pixel[522];
      node1482_l = node1474_r & ~pixel[522];
      node1483_r = node1482_l & pixel[496];
      node1483_l = node1482_l & ~pixel[496];
      node1484 = node1483_l;
      node1485 = node1483_r;
      node1486_r = node1482_r & pixel[624];
      node1486_l = node1482_r & ~pixel[624];
      node1487 = node1486_l;
      node1488 = node1486_r;
      node1489_r = node1473_r & pixel[434];
      node1489_l = node1473_r & ~pixel[434];
      node1490_r = node1489_l & pixel[629];
      node1490_l = node1489_l & ~pixel[629];
      node1491_r = node1490_l & pixel[152];
      node1491_l = node1490_l & ~pixel[152];
      node1492 = node1491_l;
      node1493 = node1491_r;
      node1494_r = node1490_r & pixel[488];
      node1494_l = node1490_r & ~pixel[488];
      node1495 = node1494_l;
      node1496 = node1494_r;
      node1497_r = node1489_r & pixel[300];
      node1497_l = node1489_r & ~pixel[300];
      node1498_r = node1497_l & pixel[346];
      node1498_l = node1497_l & ~pixel[346];
      node1499 = node1498_l;
      node1500 = node1498_r;
      node1501_r = node1497_r & pixel[439];
      node1501_l = node1497_r & ~pixel[439];
      node1502 = node1501_l;
      node1503 = node1501_r;
      node1504_r = node1472_r & pixel[428];
      node1504_l = node1472_r & ~pixel[428];
      node1505_r = node1504_l & pixel[291];
      node1505_l = node1504_l & ~pixel[291];
      node1506_r = node1505_l & pixel[513];
      node1506_l = node1505_l & ~pixel[513];
      node1507_r = node1506_l & pixel[544];
      node1507_l = node1506_l & ~pixel[544];
      node1508 = node1507_l;
      node1509 = node1507_r;
      node1510_r = node1506_r & pixel[293];
      node1510_l = node1506_r & ~pixel[293];
      node1511 = node1510_l;
      node1512 = node1510_r;
      node1513_r = node1505_r & pixel[439];
      node1513_l = node1505_r & ~pixel[439];
      node1514_r = node1513_l & pixel[376];
      node1514_l = node1513_l & ~pixel[376];
      node1515 = node1514_l;
      node1516 = node1514_r;
      node1517_r = node1513_r & pixel[623];
      node1517_l = node1513_r & ~pixel[623];
      node1518 = node1517_l;
      node1519 = node1517_r;
      node1520_r = node1504_r & pixel[625];
      node1520_l = node1504_r & ~pixel[625];
      node1521_r = node1520_l & pixel[239];
      node1521_l = node1520_l & ~pixel[239];
      node1522_r = node1521_l & pixel[542];
      node1522_l = node1521_l & ~pixel[542];
      node1523 = node1522_l;
      node1524 = node1522_r;
      node1525_r = node1521_r & pixel[182];
      node1525_l = node1521_r & ~pixel[182];
      node1526 = node1525_l;
      node1527 = node1525_r;
      node1528_r = node1520_r & pixel[413];
      node1528_l = node1520_r & ~pixel[413];
      node1529_r = node1528_l & pixel[658];
      node1529_l = node1528_l & ~pixel[658];
      node1530 = node1529_l;
      node1531 = node1529_r;
      node1532_r = node1528_r & pixel[266];
      node1532_l = node1528_r & ~pixel[266];
      node1533 = node1532_l;
      node1534 = node1532_r;
      node1535_r = node1471_r & pixel[659];
      node1535_l = node1471_r & ~pixel[659];
      node1536_r = node1535_l & pixel[441];
      node1536_l = node1535_l & ~pixel[441];
      node1537_r = node1536_l & pixel[511];
      node1537_l = node1536_l & ~pixel[511];
      node1538_r = node1537_l & pixel[692];
      node1538_l = node1537_l & ~pixel[692];
      node1539_r = node1538_l & pixel[183];
      node1539_l = node1538_l & ~pixel[183];
      node1540 = node1539_l;
      node1541 = node1539_r;
      node1542 = node1538_r;
      node1543 = node1537_r;
      node1544_r = node1536_r & pixel[496];
      node1544_l = node1536_r & ~pixel[496];
      node1545_r = node1544_l & pixel[300];
      node1545_l = node1544_l & ~pixel[300];
      node1546 = node1545_l;
      node1547 = node1545_r;
      node1548 = node1544_r;
      node1549_r = node1535_r & pixel[430];
      node1549_l = node1535_r & ~pixel[430];
      node1550_r = node1549_l & pixel[319];
      node1550_l = node1549_l & ~pixel[319];
      node1551_r = node1550_l & pixel[583];
      node1551_l = node1550_l & ~pixel[583];
      node1552_r = node1551_l & pixel[575];
      node1552_l = node1551_l & ~pixel[575];
      node1553 = node1552_l;
      node1554 = node1552_r;
      node1555 = node1551_r;
      node1556_r = node1550_r & pixel[262];
      node1556_l = node1550_r & ~pixel[262];
      node1557 = node1556_l;
      node1558_r = node1556_r & pixel[399];
      node1558_l = node1556_r & ~pixel[399];
      node1559 = node1558_l;
      node1560 = node1558_r;
      node1561_r = node1549_r & pixel[135];
      node1561_l = node1549_r & ~pixel[135];
      node1562_r = node1561_l & pixel[679];
      node1562_l = node1561_l & ~pixel[679];
      node1563_r = node1562_l & pixel[388];
      node1563_l = node1562_l & ~pixel[388];
      node1564 = node1563_l;
      node1565 = node1563_r;
      node1566 = node1562_r;
      node1567_r = node1561_r & pixel[569];
      node1567_l = node1561_r & ~pixel[569];
      node1568 = node1567_l;
      node1569 = node1567_r;
      node1570_r = node1470_r & pixel[544];
      node1570_l = node1470_r & ~pixel[544];
      node1571_r = node1570_l & pixel[484];
      node1571_l = node1570_l & ~pixel[484];
      node1572_r = node1571_l & pixel[327];
      node1572_l = node1571_l & ~pixel[327];
      node1573_r = node1572_l & pixel[297];
      node1573_l = node1572_l & ~pixel[297];
      node1574_r = node1573_l & pixel[213];
      node1574_l = node1573_l & ~pixel[213];
      node1575_r = node1574_l & pixel[513];
      node1575_l = node1574_l & ~pixel[513];
      node1576 = node1575_l;
      node1577 = node1575_r;
      node1578_r = node1574_r & pixel[147];
      node1578_l = node1574_r & ~pixel[147];
      node1579 = node1578_l;
      node1580 = node1578_r;
      node1581_r = node1573_r & pixel[514];
      node1581_l = node1573_r & ~pixel[514];
      node1582_r = node1581_l & pixel[219];
      node1582_l = node1581_l & ~pixel[219];
      node1583 = node1582_l;
      node1584 = node1582_r;
      node1585_r = node1581_r & pixel[566];
      node1585_l = node1581_r & ~pixel[566];
      node1586 = node1585_l;
      node1587 = node1585_r;
      node1588_r = node1572_r & pixel[346];
      node1588_l = node1572_r & ~pixel[346];
      node1589_r = node1588_l & pixel[594];
      node1589_l = node1588_l & ~pixel[594];
      node1590_r = node1589_l & pixel[607];
      node1590_l = node1589_l & ~pixel[607];
      node1591 = node1590_l;
      node1592 = node1590_r;
      node1593_r = node1589_r & pixel[352];
      node1593_l = node1589_r & ~pixel[352];
      node1594 = node1593_l;
      node1595 = node1593_r;
      node1596_r = node1588_r & pixel[594];
      node1596_l = node1588_r & ~pixel[594];
      node1597_r = node1596_l & pixel[412];
      node1597_l = node1596_l & ~pixel[412];
      node1598 = node1597_l;
      node1599 = node1597_r;
      node1600_r = node1596_r & pixel[348];
      node1600_l = node1596_r & ~pixel[348];
      node1601 = node1600_l;
      node1602 = node1600_r;
      node1603_r = node1571_r & pixel[377];
      node1603_l = node1571_r & ~pixel[377];
      node1604_r = node1603_l & pixel[131];
      node1604_l = node1603_l & ~pixel[131];
      node1605_r = node1604_l & pixel[628];
      node1605_l = node1604_l & ~pixel[628];
      node1606_r = node1605_l & pixel[662];
      node1606_l = node1605_l & ~pixel[662];
      node1607 = node1606_l;
      node1608 = node1606_r;
      node1609_r = node1605_r & pixel[464];
      node1609_l = node1605_r & ~pixel[464];
      node1610 = node1609_l;
      node1611 = node1609_r;
      node1612_r = node1604_r & pixel[355];
      node1612_l = node1604_r & ~pixel[355];
      node1613_r = node1612_l & pixel[513];
      node1613_l = node1612_l & ~pixel[513];
      node1614 = node1613_l;
      node1615 = node1613_r;
      node1616_r = node1612_r & pixel[467];
      node1616_l = node1612_r & ~pixel[467];
      node1617 = node1616_l;
      node1618 = node1616_r;
      node1619_r = node1603_r & pixel[345];
      node1619_l = node1603_r & ~pixel[345];
      node1620_r = node1619_l & pixel[547];
      node1620_l = node1619_l & ~pixel[547];
      node1621_r = node1620_l & pixel[320];
      node1621_l = node1620_l & ~pixel[320];
      node1622 = node1621_l;
      node1623 = node1621_r;
      node1624_r = node1620_r & pixel[679];
      node1624_l = node1620_r & ~pixel[679];
      node1625 = node1624_l;
      node1626 = node1624_r;
      node1627_r = node1619_r & pixel[273];
      node1627_l = node1619_r & ~pixel[273];
      node1628_r = node1627_l & pixel[574];
      node1628_l = node1627_l & ~pixel[574];
      node1629 = node1628_l;
      node1630 = node1628_r;
      node1631_r = node1627_r & pixel[434];
      node1631_l = node1627_r & ~pixel[434];
      node1632 = node1631_l;
      node1633 = node1631_r;
      node1634_r = node1570_r & pixel[299];
      node1634_l = node1570_r & ~pixel[299];
      node1635_r = node1634_l & pixel[429];
      node1635_l = node1634_l & ~pixel[429];
      node1636_r = node1635_l & pixel[329];
      node1636_l = node1635_l & ~pixel[329];
      node1637_r = node1636_l & pixel[346];
      node1637_l = node1636_l & ~pixel[346];
      node1638_r = node1637_l & pixel[102];
      node1638_l = node1637_l & ~pixel[102];
      node1639 = node1638_l;
      node1640 = node1638_r;
      node1641_r = node1637_r & pixel[206];
      node1641_l = node1637_r & ~pixel[206];
      node1642 = node1641_l;
      node1643 = node1641_r;
      node1644_r = node1636_r & pixel[685];
      node1644_l = node1636_r & ~pixel[685];
      node1645 = node1644_l;
      node1646 = node1644_r;
      node1647_r = node1635_r & pixel[297];
      node1647_l = node1635_r & ~pixel[297];
      node1648_r = node1647_l & pixel[191];
      node1648_l = node1647_l & ~pixel[191];
      node1649_r = node1648_l & pixel[102];
      node1649_l = node1648_l & ~pixel[102];
      node1650 = node1649_l;
      node1651 = node1649_r;
      node1652_r = node1648_r & pixel[247];
      node1652_l = node1648_r & ~pixel[247];
      node1653 = node1652_l;
      node1654 = node1652_r;
      node1655_r = node1647_r & pixel[630];
      node1655_l = node1647_r & ~pixel[630];
      node1656_r = node1655_l & pixel[156];
      node1656_l = node1655_l & ~pixel[156];
      node1657 = node1656_l;
      node1658 = node1656_r;
      node1659_r = node1655_r & pixel[359];
      node1659_l = node1655_r & ~pixel[359];
      node1660 = node1659_l;
      node1661 = node1659_r;
      node1662_r = node1634_r & pixel[348];
      node1662_l = node1634_r & ~pixel[348];
      node1663_r = node1662_l & pixel[414];
      node1663_l = node1662_l & ~pixel[414];
      node1664_r = node1663_l & pixel[183];
      node1664_l = node1663_l & ~pixel[183];
      node1665_r = node1664_l & pixel[655];
      node1665_l = node1664_l & ~pixel[655];
      node1666 = node1665_l;
      node1667 = node1665_r;
      node1668_r = node1664_r & pixel[661];
      node1668_l = node1664_r & ~pixel[661];
      node1669 = node1668_l;
      node1670 = node1668_r;
      node1671_r = node1663_r & pixel[653];
      node1671_l = node1663_r & ~pixel[653];
      node1672_r = node1671_l & pixel[688];
      node1672_l = node1671_l & ~pixel[688];
      node1673 = node1672_l;
      node1674 = node1672_r;
      node1675_r = node1671_r & pixel[350];
      node1675_l = node1671_r & ~pixel[350];
      node1676 = node1675_l;
      node1677 = node1675_r;
      node1678_r = node1662_r & pixel[358];
      node1678_l = node1662_r & ~pixel[358];
      node1679_r = node1678_l & pixel[101];
      node1679_l = node1678_l & ~pixel[101];
      node1680_r = node1679_l & pixel[628];
      node1680_l = node1679_l & ~pixel[628];
      node1681 = node1680_l;
      node1682 = node1680_r;
      node1683_r = node1679_r & pixel[180];
      node1683_l = node1679_r & ~pixel[180];
      node1684 = node1683_l;
      node1685 = node1683_r;
      node1686_r = node1678_r & pixel[274];
      node1686_l = node1678_r & ~pixel[274];
      node1687_r = node1686_l & pixel[636];
      node1687_l = node1686_l & ~pixel[636];
      node1688 = node1687_l;
      node1689 = node1687_r;
      node1690_r = node1686_r & pixel[431];
      node1690_l = node1686_r & ~pixel[431];
      node1691 = node1690_l;
      node1692 = node1690_r;
      result0 = node32 | node52 | node60 | node67 | node84 | node108 | node141 | node152 | node160 | node163 | node170 | node173 | node174 | node176 | node177 | node206 | node237 | node271 | node284 | node299 | node308 | node324 | node384 | node395 | node407 | node411 | node422 | node426 | node433 | node439 | node440 | node449 | node454 | node461 | node485 | node488 | node491 | node492 | node502 | node505 | node508 | node514 | node517 | node518 | node521 | node522 | node524 | node525 | node536 | node544 | node551 | node554 | node570 | node587 | node592 | node596 | node600 | node603 | node610 | node611 | node618 | node622 | node625 | node628 | node633 | node634 | node640 | node641 | node646 | node654 | node656 | node659 | node671 | node683 | node686 | node696 | node705 | node709 | node714 | node716 | node718 | node721 | node725 | node728 | node729 | node747 | node763 | node772 | node801 | node810 | node826 | node832 | node889 | node948 | node1012 | node1336 | node1565 | node1587 | node1610 | node1632 | node1661 | node1677 | node1692;
      result1 = node368 | node843 | node844 | node861 | node865 | node878 | node900 | node915 | node919 | node978 | node1312 | node1325 | node1436 | node1451 | node1553 | node1640;
      result2 = node26 | node33 | node44 | node48 | node49 | node56 | node63 | node64 | node92 | node96 | node107 | node119 | node120 | node122 | node129 | node137 | node138 | node140 | node144 | node159 | node169 | node181 | node192 | node208 | node232 | node245 | node248 | node267 | node287 | node296 | node302 | node307 | node309 | node345 | node353 | node355 | node360 | node361 | node364 | node401 | node402 | node415 | node418 | node429 | node457 | node510 | node533 | node648 | node670 | node673 | node674 | node744 | node760 | node769 | node771 | node783 | node791 | node798 | node802 | node829 | node847 | node875 | node884 | node901 | node907 | node911 | node924 | node929 | node959 | node964 | node967 | node974 | node981 | node1013 | node1022 | node1026 | node1027 | node1029 | node1038 | node1054 | node1060 | node1065 | node1068 | node1073 | node1076 | node1094 | node1100 | node1103 | node1106 | node1107 | node1196 | node1198 | node1202 | node1213 | node1226 | node1227 | node1230 | node1232 | node1236 | node1253 | node1261 | node1280 | node1326 | node1437 | node1439 | node1462 | node1466 | node1468 | node1478 | node1485 | node1493 | node1540 | node1541 | node1543 | node1554 | node1555 | node1566 | node1594 | node1607 | node1617 | node1625 | node1639 | node1658 | node1666 | node1669 | node1670 | node1676 | node1681 | node1685;
      result3 = node11 | node21 | node36 | node41 | node45 | node57 | node59 | node66 | node80 | node91 | node127 | node168 | node201 | node202 | node205 | node217 | node223 | node229 | node233 | node239 | node244 | node247 | node252 | node254 | node380 | node392 | node468 | node471 | node571 | node577 | node581 | node584 | node588 | node593 | node595 | node619 | node636 | node662 | node684 | node687 | node768 | node874 | node923 | node930 | node932 | node933 | node937 | node938 | node945 | node962 | node966 | node982 | node998 | node1020 | node1023 | node1034 | node1037 | node1050 | node1051 | node1053 | node1058 | node1061 | node1069 | node1072 | node1085 | node1087 | node1091 | node1102 | node1108 | node1132 | node1135 | node1167 | node1185 | node1205 | node1210 | node1214 | node1239 | node1279 | node1287 | node1343 | node1373 | node1376 | node1382 | node1383 | node1453 | node1508 | node1509 | node1519 | node1530 | node1557 | node1583 | node1591 | node1595 | node1602 | node1622 | node1626 | node1689;
      result4 = node20 | node28 | node83 | node112 | node153 | node156 | node209 | node276 | node279 | node310 | node319 | node333 | node336 | node346 | node352 | node369 | node398 | node414 | node463 | node478 | node483 | node484 | node537 | node543 | node563 | node615 | node649 | node693 | node708 | node715 | node730 | node741 | node752 | node759 | node778 | node784 | node786 | node799 | node807 | node823 | node881 | node885 | node892 | node916 | node958 | node975 | node987 | node991 | node995 | node1010 | node1084 | node1099 | node1113 | node1120 | node1131 | node1143 | node1146 | node1156 | node1246 | node1249 | node1257 | node1266 | node1274 | node1296 | node1297 | node1313 | node1319 | node1348 | node1388 | node1392 | node1397 | node1523 | node1524 | node1526 | node1533 | node1548 | node1608 | node1657;
      result5 = node10 | node14 | node29 | node35 | node42 | node99 | node111 | node115 | node123 | node126 | node147 | node198 | node199 | node213 | node214 | node220 | node224 | node230 | node236 | node240 | node251 | node255 | node263 | node270 | node327 | node376 | node377 | node379 | node383 | node387 | node391 | node408 | node423 | node430 | node447 | node469 | node472 | node475 | node476 | node489 | node567 | node580 | node585 | node599 | node602 | node612 | node616 | node627 | node637 | node661 | node694 | node850 | node853 | node858 | node859 | node882 | node888 | node893 | node904 | node942 | node950 | node1005 | node1041 | node1044 | node1117 | node1124 | node1129 | node1137 | node1152 | node1165 | node1172 | node1179 | node1188 | node1269 | node1277 | node1284 | node1328 | node1332 | node1335 | node1358 | node1401 | node1411 | node1419 | node1446 | node1477 | node1481 | node1488 | node1492 | node1495 | node1560 | node1569 | node1576 | node1577 | node1579 | node1580 | node1584 | node1599 | node1611 | node1614 | node1629 | node1642 | node1643 | node1653;
      result6 = node25 | node51 | node162 | node184 | node216 | node264 | node266 | node280 | node292 | node293 | node295 | node300 | node303 | node323 | node326 | node356 | node363 | node366 | node386 | node479 | node504 | node515 | node530 | node534 | node540 | node542 | node556 | node564 | node566 | node572 | node578 | node624 | node681 | node682 | node697 | node699 | node701 | node702 | node737 | node738 | node745 | node748 | node762 | node780 | node811 | node817 | node822 | node854 | node877 | node894 | node903 | node908 | node910 | node971 | node972 | node988 | node990 | node1003 | node1019 | node1030 | node1114 | node1121 | node1144 | node1148 | node1151 | node1159 | node1181 | node1199 | node1203 | node1238 | node1240 | node1247 | node1250 | node1256 | node1267 | node1298 | node1305 | node1309 | node1310 | node1320 | node1420 | node1422 | node1423 | node1426 | node1427 | node1428 | node1432 | node1434 | node1440 | node1447 | node1448 | node1452 | node1457 | node1458 | node1463 | node1464 | node1469 | node1487 | node1496 | node1500 | node1534 | node1546 | node1568 | node1615 | node1630 | node1645 | node1650 | node1651 | node1654 | node1673 | node1684 | node1688;
      result7 = node13 | node17 | node18 | node73 | node74 | node76 | node77 | node81 | node88 | node105 | node277 | node316 | node317 | node339 | node349 | node394 | node399 | node410 | node442 | node446 | node501 | node509 | node550 | node553 | node559 | node644 | node651 | node657 | node675 | node753 | node755 | node794 | node795 | node815 | node818 | node833 | node846 | node979 | node1195 | node1211 | node1262 | node1351 | node1361 | node1364 | node1372 | node1375 | node1379 | node1389 | node1396;
      result8 = node130 | node148 | node182 | node188 | node189 | node191 | node221 | node272 | node425 | node432 | node450 | node458 | node462 | node531 | node558 | node740 | node770 | node787 | node830 | node862 | node866 | node868 | node869 | node918 | node936 | node943 | node946 | node951 | node994 | node997 | node1002 | node1035 | node1042 | node1045 | node1057 | node1066 | node1075 | node1088 | node1092 | node1095 | node1123 | node1128 | node1136 | node1155 | node1158 | node1168 | node1171 | node1175 | node1180 | node1187 | node1206 | node1217 | node1218 | node1220 | node1221 | node1229 | node1233 | node1254 | node1263 | node1270 | node1273 | node1283 | node1286 | node1302 | node1304 | node1316 | node1317 | node1329 | node1333 | node1341 | node1344 | node1360 | node1405 | node1408 | node1412 | node1431 | node1456 | node1480 | node1484 | node1499 | node1502 | node1503 | node1511 | node1512 | node1515 | node1516 | node1518 | node1531 | node1542 | node1559 | node1564 | node1586 | node1592 | node1598 | node1618 | node1623 | node1633 | node1646 | node1660 | node1667 | node1682 | node1691;
      result9 = node89 | node95 | node98 | node104 | node114 | node145 | node155 | node185 | node283 | node286 | node320 | node330 | node332 | node337 | node340 | node348 | node417 | node443 | node455 | node643 | node676 | node706 | node720 | node724 | node756 | node779 | node792 | node808 | node814 | node825 | node851 | node922 | node961 | node1006 | node1009 | node1116 | node1147 | node1164 | node1174 | node1184 | node1301 | node1340 | node1347 | node1350 | node1357 | node1365 | node1367 | node1368 | node1380 | node1391 | node1394 | node1402 | node1404 | node1409 | node1527 | node1547 | node1601 | node1674;

      tree_6 = {result9, result8, result7, result6, result5, result4, result3, result2, result1, result0};
    end
  endfunction

  function [9:0] tree_7;
    input [783:0] pixel;

    reg node0_r;
    reg node0_l;
    reg node1_r;
    reg node1_l;
    reg node2_r;
    reg node2_l;
    reg node3_r;
    reg node3_l;
    reg node4_r;
    reg node4_l;
    reg node5_r;
    reg node5_l;
    reg node6_r;
    reg node6_l;
    reg node7_r;
    reg node7_l;
    reg node8_r;
    reg node8_l;
    reg node9_r;
    reg node9_l;
    reg node10;
    reg node11;
    reg node12_r;
    reg node12_l;
    reg node13;
    reg node14;
    reg node15_r;
    reg node15_l;
    reg node16_r;
    reg node16_l;
    reg node17;
    reg node18;
    reg node19_r;
    reg node19_l;
    reg node20;
    reg node21;
    reg node22_r;
    reg node22_l;
    reg node23_r;
    reg node23_l;
    reg node24_r;
    reg node24_l;
    reg node25;
    reg node26;
    reg node27_r;
    reg node27_l;
    reg node28;
    reg node29;
    reg node30_r;
    reg node30_l;
    reg node31_r;
    reg node31_l;
    reg node32;
    reg node33;
    reg node34_r;
    reg node34_l;
    reg node35;
    reg node36;
    reg node37_r;
    reg node37_l;
    reg node38_r;
    reg node38_l;
    reg node39_r;
    reg node39_l;
    reg node40_r;
    reg node40_l;
    reg node41;
    reg node42;
    reg node43_r;
    reg node43_l;
    reg node44;
    reg node45;
    reg node46_r;
    reg node46_l;
    reg node47_r;
    reg node47_l;
    reg node48;
    reg node49;
    reg node50_r;
    reg node50_l;
    reg node51;
    reg node52;
    reg node53_r;
    reg node53_l;
    reg node54_r;
    reg node54_l;
    reg node55_r;
    reg node55_l;
    reg node56;
    reg node57;
    reg node58;
    reg node59_r;
    reg node59_l;
    reg node60;
    reg node61_r;
    reg node61_l;
    reg node62;
    reg node63;
    reg node64_r;
    reg node64_l;
    reg node65_r;
    reg node65_l;
    reg node66_r;
    reg node66_l;
    reg node67_r;
    reg node67_l;
    reg node68_r;
    reg node68_l;
    reg node69;
    reg node70;
    reg node71_r;
    reg node71_l;
    reg node72;
    reg node73;
    reg node74_r;
    reg node74_l;
    reg node75;
    reg node76_r;
    reg node76_l;
    reg node77;
    reg node78;
    reg node79_r;
    reg node79_l;
    reg node80_r;
    reg node80_l;
    reg node81_r;
    reg node81_l;
    reg node82;
    reg node83;
    reg node84_r;
    reg node84_l;
    reg node85;
    reg node86;
    reg node87_r;
    reg node87_l;
    reg node88_r;
    reg node88_l;
    reg node89;
    reg node90;
    reg node91_r;
    reg node91_l;
    reg node92;
    reg node93;
    reg node94_r;
    reg node94_l;
    reg node95_r;
    reg node95_l;
    reg node96_r;
    reg node96_l;
    reg node97_r;
    reg node97_l;
    reg node98;
    reg node99;
    reg node100_r;
    reg node100_l;
    reg node101;
    reg node102;
    reg node103_r;
    reg node103_l;
    reg node104_r;
    reg node104_l;
    reg node105;
    reg node106;
    reg node107_r;
    reg node107_l;
    reg node108;
    reg node109;
    reg node110_r;
    reg node110_l;
    reg node111_r;
    reg node111_l;
    reg node112_r;
    reg node112_l;
    reg node113;
    reg node114;
    reg node115_r;
    reg node115_l;
    reg node116;
    reg node117;
    reg node118_r;
    reg node118_l;
    reg node119_r;
    reg node119_l;
    reg node120;
    reg node121;
    reg node122_r;
    reg node122_l;
    reg node123;
    reg node124;
    reg node125_r;
    reg node125_l;
    reg node126_r;
    reg node126_l;
    reg node127_r;
    reg node127_l;
    reg node128_r;
    reg node128_l;
    reg node129_r;
    reg node129_l;
    reg node130_r;
    reg node130_l;
    reg node131;
    reg node132;
    reg node133_r;
    reg node133_l;
    reg node134;
    reg node135;
    reg node136_r;
    reg node136_l;
    reg node137_r;
    reg node137_l;
    reg node138;
    reg node139;
    reg node140_r;
    reg node140_l;
    reg node141;
    reg node142;
    reg node143_r;
    reg node143_l;
    reg node144_r;
    reg node144_l;
    reg node145_r;
    reg node145_l;
    reg node146;
    reg node147;
    reg node148_r;
    reg node148_l;
    reg node149;
    reg node150;
    reg node151_r;
    reg node151_l;
    reg node152_r;
    reg node152_l;
    reg node153;
    reg node154;
    reg node155_r;
    reg node155_l;
    reg node156;
    reg node157;
    reg node158_r;
    reg node158_l;
    reg node159_r;
    reg node159_l;
    reg node160_r;
    reg node160_l;
    reg node161_r;
    reg node161_l;
    reg node162;
    reg node163;
    reg node164_r;
    reg node164_l;
    reg node165;
    reg node166;
    reg node167_r;
    reg node167_l;
    reg node168_r;
    reg node168_l;
    reg node169;
    reg node170;
    reg node171_r;
    reg node171_l;
    reg node172;
    reg node173;
    reg node174_r;
    reg node174_l;
    reg node175_r;
    reg node175_l;
    reg node176_r;
    reg node176_l;
    reg node177;
    reg node178;
    reg node179_r;
    reg node179_l;
    reg node180;
    reg node181;
    reg node182_r;
    reg node182_l;
    reg node183_r;
    reg node183_l;
    reg node184;
    reg node185;
    reg node186_r;
    reg node186_l;
    reg node187;
    reg node188;
    reg node189_r;
    reg node189_l;
    reg node190_r;
    reg node190_l;
    reg node191;
    reg node192_r;
    reg node192_l;
    reg node193_r;
    reg node193_l;
    reg node194;
    reg node195_r;
    reg node195_l;
    reg node196;
    reg node197;
    reg node198;
    reg node199_r;
    reg node199_l;
    reg node200_r;
    reg node200_l;
    reg node201_r;
    reg node201_l;
    reg node202;
    reg node203_r;
    reg node203_l;
    reg node204;
    reg node205;
    reg node206_r;
    reg node206_l;
    reg node207;
    reg node208;
    reg node209_r;
    reg node209_l;
    reg node210_r;
    reg node210_l;
    reg node211_r;
    reg node211_l;
    reg node212;
    reg node213;
    reg node214_r;
    reg node214_l;
    reg node215;
    reg node216;
    reg node217;
    reg node218_r;
    reg node218_l;
    reg node219_r;
    reg node219_l;
    reg node220_r;
    reg node220_l;
    reg node221_r;
    reg node221_l;
    reg node222_r;
    reg node222_l;
    reg node223_r;
    reg node223_l;
    reg node224_r;
    reg node224_l;
    reg node225;
    reg node226;
    reg node227_r;
    reg node227_l;
    reg node228;
    reg node229;
    reg node230_r;
    reg node230_l;
    reg node231_r;
    reg node231_l;
    reg node232;
    reg node233;
    reg node234_r;
    reg node234_l;
    reg node235;
    reg node236;
    reg node237_r;
    reg node237_l;
    reg node238_r;
    reg node238_l;
    reg node239_r;
    reg node239_l;
    reg node240;
    reg node241;
    reg node242_r;
    reg node242_l;
    reg node243;
    reg node244;
    reg node245_r;
    reg node245_l;
    reg node246_r;
    reg node246_l;
    reg node247;
    reg node248;
    reg node249;
    reg node250_r;
    reg node250_l;
    reg node251_r;
    reg node251_l;
    reg node252_r;
    reg node252_l;
    reg node253_r;
    reg node253_l;
    reg node254;
    reg node255;
    reg node256;
    reg node257_r;
    reg node257_l;
    reg node258_r;
    reg node258_l;
    reg node259;
    reg node260;
    reg node261;
    reg node262_r;
    reg node262_l;
    reg node263;
    reg node264_r;
    reg node264_l;
    reg node265;
    reg node266;
    reg node267_r;
    reg node267_l;
    reg node268_r;
    reg node268_l;
    reg node269_r;
    reg node269_l;
    reg node270;
    reg node271_r;
    reg node271_l;
    reg node272_r;
    reg node272_l;
    reg node273;
    reg node274;
    reg node275_r;
    reg node275_l;
    reg node276;
    reg node277;
    reg node278_r;
    reg node278_l;
    reg node279_r;
    reg node279_l;
    reg node280;
    reg node281_r;
    reg node281_l;
    reg node282;
    reg node283;
    reg node284_r;
    reg node284_l;
    reg node285_r;
    reg node285_l;
    reg node286;
    reg node287;
    reg node288;
    reg node289_r;
    reg node289_l;
    reg node290_r;
    reg node290_l;
    reg node291_r;
    reg node291_l;
    reg node292_r;
    reg node292_l;
    reg node293;
    reg node294;
    reg node295_r;
    reg node295_l;
    reg node296;
    reg node297;
    reg node298_r;
    reg node298_l;
    reg node299;
    reg node300_r;
    reg node300_l;
    reg node301;
    reg node302;
    reg node303_r;
    reg node303_l;
    reg node304_r;
    reg node304_l;
    reg node305;
    reg node306_r;
    reg node306_l;
    reg node307;
    reg node308;
    reg node309_r;
    reg node309_l;
    reg node310;
    reg node311;
    reg node312_r;
    reg node312_l;
    reg node313_r;
    reg node313_l;
    reg node314_r;
    reg node314_l;
    reg node315_r;
    reg node315_l;
    reg node316_r;
    reg node316_l;
    reg node317_r;
    reg node317_l;
    reg node318;
    reg node319;
    reg node320;
    reg node321_r;
    reg node321_l;
    reg node322_r;
    reg node322_l;
    reg node323;
    reg node324;
    reg node325;
    reg node326_r;
    reg node326_l;
    reg node327_r;
    reg node327_l;
    reg node328_r;
    reg node328_l;
    reg node329;
    reg node330;
    reg node331;
    reg node332_r;
    reg node332_l;
    reg node333;
    reg node334_r;
    reg node334_l;
    reg node335;
    reg node336;
    reg node337_r;
    reg node337_l;
    reg node338_r;
    reg node338_l;
    reg node339_r;
    reg node339_l;
    reg node340_r;
    reg node340_l;
    reg node341;
    reg node342;
    reg node343_r;
    reg node343_l;
    reg node344;
    reg node345;
    reg node346_r;
    reg node346_l;
    reg node347;
    reg node348_r;
    reg node348_l;
    reg node349;
    reg node350;
    reg node351_r;
    reg node351_l;
    reg node352;
    reg node353_r;
    reg node353_l;
    reg node354_r;
    reg node354_l;
    reg node355;
    reg node356;
    reg node357_r;
    reg node357_l;
    reg node358;
    reg node359;
    reg node360_r;
    reg node360_l;
    reg node361_r;
    reg node361_l;
    reg node362_r;
    reg node362_l;
    reg node363_r;
    reg node363_l;
    reg node364_r;
    reg node364_l;
    reg node365;
    reg node366;
    reg node367;
    reg node368_r;
    reg node368_l;
    reg node369;
    reg node370;
    reg node371_r;
    reg node371_l;
    reg node372_r;
    reg node372_l;
    reg node373;
    reg node374;
    reg node375_r;
    reg node375_l;
    reg node376_r;
    reg node376_l;
    reg node377;
    reg node378;
    reg node379_r;
    reg node379_l;
    reg node380;
    reg node381;
    reg node382_r;
    reg node382_l;
    reg node383_r;
    reg node383_l;
    reg node384;
    reg node385_r;
    reg node385_l;
    reg node386;
    reg node387;
    reg node388_r;
    reg node388_l;
    reg node389_r;
    reg node389_l;
    reg node390;
    reg node391_r;
    reg node391_l;
    reg node392;
    reg node393;
    reg node394_r;
    reg node394_l;
    reg node395;
    reg node396;
    reg node397_r;
    reg node397_l;
    reg node398_r;
    reg node398_l;
    reg node399_r;
    reg node399_l;
    reg node400_r;
    reg node400_l;
    reg node401_r;
    reg node401_l;
    reg node402_r;
    reg node402_l;
    reg node403_r;
    reg node403_l;
    reg node404_r;
    reg node404_l;
    reg node405;
    reg node406;
    reg node407_r;
    reg node407_l;
    reg node408;
    reg node409;
    reg node410_r;
    reg node410_l;
    reg node411_r;
    reg node411_l;
    reg node412;
    reg node413;
    reg node414_r;
    reg node414_l;
    reg node415;
    reg node416;
    reg node417_r;
    reg node417_l;
    reg node418_r;
    reg node418_l;
    reg node419_r;
    reg node419_l;
    reg node420;
    reg node421;
    reg node422_r;
    reg node422_l;
    reg node423;
    reg node424;
    reg node425_r;
    reg node425_l;
    reg node426_r;
    reg node426_l;
    reg node427;
    reg node428;
    reg node429_r;
    reg node429_l;
    reg node430;
    reg node431;
    reg node432_r;
    reg node432_l;
    reg node433_r;
    reg node433_l;
    reg node434_r;
    reg node434_l;
    reg node435_r;
    reg node435_l;
    reg node436;
    reg node437;
    reg node438_r;
    reg node438_l;
    reg node439;
    reg node440;
    reg node441_r;
    reg node441_l;
    reg node442_r;
    reg node442_l;
    reg node443;
    reg node444;
    reg node445_r;
    reg node445_l;
    reg node446;
    reg node447;
    reg node448_r;
    reg node448_l;
    reg node449_r;
    reg node449_l;
    reg node450_r;
    reg node450_l;
    reg node451;
    reg node452;
    reg node453;
    reg node454_r;
    reg node454_l;
    reg node455;
    reg node456;
    reg node457_r;
    reg node457_l;
    reg node458_r;
    reg node458_l;
    reg node459_r;
    reg node459_l;
    reg node460_r;
    reg node460_l;
    reg node461_r;
    reg node461_l;
    reg node462;
    reg node463;
    reg node464_r;
    reg node464_l;
    reg node465;
    reg node466;
    reg node467_r;
    reg node467_l;
    reg node468_r;
    reg node468_l;
    reg node469;
    reg node470;
    reg node471_r;
    reg node471_l;
    reg node472;
    reg node473;
    reg node474_r;
    reg node474_l;
    reg node475_r;
    reg node475_l;
    reg node476_r;
    reg node476_l;
    reg node477;
    reg node478;
    reg node479_r;
    reg node479_l;
    reg node480;
    reg node481;
    reg node482_r;
    reg node482_l;
    reg node483_r;
    reg node483_l;
    reg node484;
    reg node485;
    reg node486_r;
    reg node486_l;
    reg node487;
    reg node488;
    reg node489_r;
    reg node489_l;
    reg node490_r;
    reg node490_l;
    reg node491_r;
    reg node491_l;
    reg node492_r;
    reg node492_l;
    reg node493;
    reg node494;
    reg node495_r;
    reg node495_l;
    reg node496;
    reg node497;
    reg node498_r;
    reg node498_l;
    reg node499_r;
    reg node499_l;
    reg node500;
    reg node501;
    reg node502_r;
    reg node502_l;
    reg node503;
    reg node504;
    reg node505_r;
    reg node505_l;
    reg node506_r;
    reg node506_l;
    reg node507_r;
    reg node507_l;
    reg node508;
    reg node509;
    reg node510_r;
    reg node510_l;
    reg node511;
    reg node512;
    reg node513_r;
    reg node513_l;
    reg node514_r;
    reg node514_l;
    reg node515;
    reg node516;
    reg node517;
    reg node518_r;
    reg node518_l;
    reg node519_r;
    reg node519_l;
    reg node520_r;
    reg node520_l;
    reg node521_r;
    reg node521_l;
    reg node522_r;
    reg node522_l;
    reg node523_r;
    reg node523_l;
    reg node524;
    reg node525;
    reg node526_r;
    reg node526_l;
    reg node527;
    reg node528;
    reg node529_r;
    reg node529_l;
    reg node530_r;
    reg node530_l;
    reg node531;
    reg node532;
    reg node533_r;
    reg node533_l;
    reg node534;
    reg node535;
    reg node536_r;
    reg node536_l;
    reg node537_r;
    reg node537_l;
    reg node538_r;
    reg node538_l;
    reg node539;
    reg node540;
    reg node541;
    reg node542_r;
    reg node542_l;
    reg node543_r;
    reg node543_l;
    reg node544;
    reg node545;
    reg node546_r;
    reg node546_l;
    reg node547;
    reg node548;
    reg node549_r;
    reg node549_l;
    reg node550_r;
    reg node550_l;
    reg node551_r;
    reg node551_l;
    reg node552_r;
    reg node552_l;
    reg node553;
    reg node554;
    reg node555_r;
    reg node555_l;
    reg node556;
    reg node557;
    reg node558_r;
    reg node558_l;
    reg node559_r;
    reg node559_l;
    reg node560;
    reg node561;
    reg node562_r;
    reg node562_l;
    reg node563;
    reg node564;
    reg node565_r;
    reg node565_l;
    reg node566_r;
    reg node566_l;
    reg node567_r;
    reg node567_l;
    reg node568;
    reg node569;
    reg node570_r;
    reg node570_l;
    reg node571;
    reg node572;
    reg node573_r;
    reg node573_l;
    reg node574_r;
    reg node574_l;
    reg node575;
    reg node576;
    reg node577_r;
    reg node577_l;
    reg node578;
    reg node579;
    reg node580_r;
    reg node580_l;
    reg node581_r;
    reg node581_l;
    reg node582_r;
    reg node582_l;
    reg node583_r;
    reg node583_l;
    reg node584_r;
    reg node584_l;
    reg node585;
    reg node586;
    reg node587_r;
    reg node587_l;
    reg node588;
    reg node589;
    reg node590_r;
    reg node590_l;
    reg node591_r;
    reg node591_l;
    reg node592;
    reg node593;
    reg node594_r;
    reg node594_l;
    reg node595;
    reg node596;
    reg node597_r;
    reg node597_l;
    reg node598_r;
    reg node598_l;
    reg node599_r;
    reg node599_l;
    reg node600;
    reg node601;
    reg node602_r;
    reg node602_l;
    reg node603;
    reg node604;
    reg node605_r;
    reg node605_l;
    reg node606_r;
    reg node606_l;
    reg node607;
    reg node608;
    reg node609_r;
    reg node609_l;
    reg node610;
    reg node611;
    reg node612_r;
    reg node612_l;
    reg node613_r;
    reg node613_l;
    reg node614_r;
    reg node614_l;
    reg node615_r;
    reg node615_l;
    reg node616;
    reg node617;
    reg node618_r;
    reg node618_l;
    reg node619;
    reg node620;
    reg node621_r;
    reg node621_l;
    reg node622_r;
    reg node622_l;
    reg node623;
    reg node624;
    reg node625_r;
    reg node625_l;
    reg node626;
    reg node627;
    reg node628_r;
    reg node628_l;
    reg node629_r;
    reg node629_l;
    reg node630_r;
    reg node630_l;
    reg node631;
    reg node632;
    reg node633;
    reg node634_r;
    reg node634_l;
    reg node635_r;
    reg node635_l;
    reg node636;
    reg node637;
    reg node638_r;
    reg node638_l;
    reg node639;
    reg node640;
    reg node641_r;
    reg node641_l;
    reg node642_r;
    reg node642_l;
    reg node643_r;
    reg node643_l;
    reg node644_r;
    reg node644_l;
    reg node645_r;
    reg node645_l;
    reg node646_r;
    reg node646_l;
    reg node647_r;
    reg node647_l;
    reg node648;
    reg node649;
    reg node650_r;
    reg node650_l;
    reg node651;
    reg node652;
    reg node653_r;
    reg node653_l;
    reg node654_r;
    reg node654_l;
    reg node655;
    reg node656;
    reg node657;
    reg node658_r;
    reg node658_l;
    reg node659_r;
    reg node659_l;
    reg node660_r;
    reg node660_l;
    reg node661;
    reg node662;
    reg node663_r;
    reg node663_l;
    reg node664;
    reg node665;
    reg node666_r;
    reg node666_l;
    reg node667_r;
    reg node667_l;
    reg node668;
    reg node669;
    reg node670_r;
    reg node670_l;
    reg node671;
    reg node672;
    reg node673_r;
    reg node673_l;
    reg node674_r;
    reg node674_l;
    reg node675_r;
    reg node675_l;
    reg node676_r;
    reg node676_l;
    reg node677;
    reg node678;
    reg node679_r;
    reg node679_l;
    reg node680;
    reg node681;
    reg node682_r;
    reg node682_l;
    reg node683_r;
    reg node683_l;
    reg node684;
    reg node685;
    reg node686_r;
    reg node686_l;
    reg node687;
    reg node688;
    reg node689_r;
    reg node689_l;
    reg node690_r;
    reg node690_l;
    reg node691_r;
    reg node691_l;
    reg node692;
    reg node693;
    reg node694_r;
    reg node694_l;
    reg node695;
    reg node696;
    reg node697_r;
    reg node697_l;
    reg node698_r;
    reg node698_l;
    reg node699;
    reg node700;
    reg node701_r;
    reg node701_l;
    reg node702;
    reg node703;
    reg node704_r;
    reg node704_l;
    reg node705_r;
    reg node705_l;
    reg node706_r;
    reg node706_l;
    reg node707_r;
    reg node707_l;
    reg node708_r;
    reg node708_l;
    reg node709;
    reg node710;
    reg node711_r;
    reg node711_l;
    reg node712;
    reg node713;
    reg node714_r;
    reg node714_l;
    reg node715_r;
    reg node715_l;
    reg node716;
    reg node717;
    reg node718_r;
    reg node718_l;
    reg node719;
    reg node720;
    reg node721_r;
    reg node721_l;
    reg node722_r;
    reg node722_l;
    reg node723_r;
    reg node723_l;
    reg node724;
    reg node725;
    reg node726;
    reg node727_r;
    reg node727_l;
    reg node728_r;
    reg node728_l;
    reg node729;
    reg node730;
    reg node731_r;
    reg node731_l;
    reg node732;
    reg node733;
    reg node734_r;
    reg node734_l;
    reg node735_r;
    reg node735_l;
    reg node736_r;
    reg node736_l;
    reg node737_r;
    reg node737_l;
    reg node738;
    reg node739;
    reg node740_r;
    reg node740_l;
    reg node741;
    reg node742;
    reg node743_r;
    reg node743_l;
    reg node744_r;
    reg node744_l;
    reg node745;
    reg node746;
    reg node747_r;
    reg node747_l;
    reg node748;
    reg node749;
    reg node750_r;
    reg node750_l;
    reg node751;
    reg node752_r;
    reg node752_l;
    reg node753_r;
    reg node753_l;
    reg node754;
    reg node755;
    reg node756_r;
    reg node756_l;
    reg node757;
    reg node758;
    reg node759_r;
    reg node759_l;
    reg node760_r;
    reg node760_l;
    reg node761_r;
    reg node761_l;
    reg node762_r;
    reg node762_l;
    reg node763_r;
    reg node763_l;
    reg node764_r;
    reg node764_l;
    reg node765;
    reg node766;
    reg node767_r;
    reg node767_l;
    reg node768;
    reg node769;
    reg node770_r;
    reg node770_l;
    reg node771_r;
    reg node771_l;
    reg node772;
    reg node773;
    reg node774_r;
    reg node774_l;
    reg node775;
    reg node776;
    reg node777_r;
    reg node777_l;
    reg node778_r;
    reg node778_l;
    reg node779_r;
    reg node779_l;
    reg node780;
    reg node781;
    reg node782_r;
    reg node782_l;
    reg node783;
    reg node784;
    reg node785_r;
    reg node785_l;
    reg node786_r;
    reg node786_l;
    reg node787;
    reg node788;
    reg node789_r;
    reg node789_l;
    reg node790;
    reg node791;
    reg node792_r;
    reg node792_l;
    reg node793_r;
    reg node793_l;
    reg node794_r;
    reg node794_l;
    reg node795_r;
    reg node795_l;
    reg node796;
    reg node797;
    reg node798_r;
    reg node798_l;
    reg node799;
    reg node800;
    reg node801_r;
    reg node801_l;
    reg node802_r;
    reg node802_l;
    reg node803;
    reg node804;
    reg node805_r;
    reg node805_l;
    reg node806;
    reg node807;
    reg node808_r;
    reg node808_l;
    reg node809_r;
    reg node809_l;
    reg node810_r;
    reg node810_l;
    reg node811;
    reg node812;
    reg node813_r;
    reg node813_l;
    reg node814;
    reg node815;
    reg node816_r;
    reg node816_l;
    reg node817_r;
    reg node817_l;
    reg node818;
    reg node819;
    reg node820_r;
    reg node820_l;
    reg node821;
    reg node822;
    reg node823_r;
    reg node823_l;
    reg node824_r;
    reg node824_l;
    reg node825_r;
    reg node825_l;
    reg node826_r;
    reg node826_l;
    reg node827_r;
    reg node827_l;
    reg node828;
    reg node829;
    reg node830_r;
    reg node830_l;
    reg node831;
    reg node832;
    reg node833_r;
    reg node833_l;
    reg node834_r;
    reg node834_l;
    reg node835;
    reg node836;
    reg node837_r;
    reg node837_l;
    reg node838;
    reg node839;
    reg node840_r;
    reg node840_l;
    reg node841_r;
    reg node841_l;
    reg node842_r;
    reg node842_l;
    reg node843;
    reg node844;
    reg node845_r;
    reg node845_l;
    reg node846;
    reg node847;
    reg node848_r;
    reg node848_l;
    reg node849_r;
    reg node849_l;
    reg node850;
    reg node851;
    reg node852_r;
    reg node852_l;
    reg node853;
    reg node854;
    reg node855_r;
    reg node855_l;
    reg node856_r;
    reg node856_l;
    reg node857_r;
    reg node857_l;
    reg node858;
    reg node859;
    reg node860_r;
    reg node860_l;
    reg node861;
    reg node862;
    reg node863;
    reg node864_r;
    reg node864_l;
    reg node865_r;
    reg node865_l;
    reg node866_r;
    reg node866_l;
    reg node867_r;
    reg node867_l;
    reg node868_r;
    reg node868_l;
    reg node869_r;
    reg node869_l;
    reg node870_r;
    reg node870_l;
    reg node871_r;
    reg node871_l;
    reg node872_r;
    reg node872_l;
    reg node873;
    reg node874;
    reg node875_r;
    reg node875_l;
    reg node876;
    reg node877;
    reg node878_r;
    reg node878_l;
    reg node879_r;
    reg node879_l;
    reg node880;
    reg node881;
    reg node882_r;
    reg node882_l;
    reg node883;
    reg node884;
    reg node885_r;
    reg node885_l;
    reg node886_r;
    reg node886_l;
    reg node887_r;
    reg node887_l;
    reg node888;
    reg node889;
    reg node890_r;
    reg node890_l;
    reg node891;
    reg node892;
    reg node893_r;
    reg node893_l;
    reg node894_r;
    reg node894_l;
    reg node895;
    reg node896;
    reg node897_r;
    reg node897_l;
    reg node898;
    reg node899;
    reg node900_r;
    reg node900_l;
    reg node901_r;
    reg node901_l;
    reg node902_r;
    reg node902_l;
    reg node903_r;
    reg node903_l;
    reg node904;
    reg node905;
    reg node906_r;
    reg node906_l;
    reg node907;
    reg node908;
    reg node909_r;
    reg node909_l;
    reg node910_r;
    reg node910_l;
    reg node911;
    reg node912;
    reg node913_r;
    reg node913_l;
    reg node914;
    reg node915;
    reg node916_r;
    reg node916_l;
    reg node917_r;
    reg node917_l;
    reg node918_r;
    reg node918_l;
    reg node919;
    reg node920;
    reg node921_r;
    reg node921_l;
    reg node922;
    reg node923;
    reg node924_r;
    reg node924_l;
    reg node925_r;
    reg node925_l;
    reg node926;
    reg node927;
    reg node928_r;
    reg node928_l;
    reg node929;
    reg node930;
    reg node931_r;
    reg node931_l;
    reg node932_r;
    reg node932_l;
    reg node933_r;
    reg node933_l;
    reg node934_r;
    reg node934_l;
    reg node935_r;
    reg node935_l;
    reg node936;
    reg node937;
    reg node938;
    reg node939_r;
    reg node939_l;
    reg node940_r;
    reg node940_l;
    reg node941;
    reg node942;
    reg node943_r;
    reg node943_l;
    reg node944;
    reg node945;
    reg node946_r;
    reg node946_l;
    reg node947_r;
    reg node947_l;
    reg node948_r;
    reg node948_l;
    reg node949;
    reg node950;
    reg node951;
    reg node952_r;
    reg node952_l;
    reg node953_r;
    reg node953_l;
    reg node954;
    reg node955;
    reg node956_r;
    reg node956_l;
    reg node957;
    reg node958;
    reg node959_r;
    reg node959_l;
    reg node960_r;
    reg node960_l;
    reg node961_r;
    reg node961_l;
    reg node962_r;
    reg node962_l;
    reg node963;
    reg node964;
    reg node965_r;
    reg node965_l;
    reg node966;
    reg node967;
    reg node968_r;
    reg node968_l;
    reg node969_r;
    reg node969_l;
    reg node970;
    reg node971;
    reg node972_r;
    reg node972_l;
    reg node973;
    reg node974;
    reg node975_r;
    reg node975_l;
    reg node976;
    reg node977_r;
    reg node977_l;
    reg node978_r;
    reg node978_l;
    reg node979;
    reg node980;
    reg node981_r;
    reg node981_l;
    reg node982;
    reg node983;
    reg node984_r;
    reg node984_l;
    reg node985_r;
    reg node985_l;
    reg node986_r;
    reg node986_l;
    reg node987_r;
    reg node987_l;
    reg node988_r;
    reg node988_l;
    reg node989_r;
    reg node989_l;
    reg node990;
    reg node991;
    reg node992_r;
    reg node992_l;
    reg node993;
    reg node994;
    reg node995_r;
    reg node995_l;
    reg node996_r;
    reg node996_l;
    reg node997;
    reg node998;
    reg node999;
    reg node1000_r;
    reg node1000_l;
    reg node1001_r;
    reg node1001_l;
    reg node1002;
    reg node1003;
    reg node1004_r;
    reg node1004_l;
    reg node1005;
    reg node1006;
    reg node1007_r;
    reg node1007_l;
    reg node1008_r;
    reg node1008_l;
    reg node1009_r;
    reg node1009_l;
    reg node1010_r;
    reg node1010_l;
    reg node1011;
    reg node1012;
    reg node1013_r;
    reg node1013_l;
    reg node1014;
    reg node1015;
    reg node1016_r;
    reg node1016_l;
    reg node1017_r;
    reg node1017_l;
    reg node1018;
    reg node1019;
    reg node1020_r;
    reg node1020_l;
    reg node1021;
    reg node1022;
    reg node1023_r;
    reg node1023_l;
    reg node1024_r;
    reg node1024_l;
    reg node1025_r;
    reg node1025_l;
    reg node1026;
    reg node1027;
    reg node1028_r;
    reg node1028_l;
    reg node1029;
    reg node1030;
    reg node1031_r;
    reg node1031_l;
    reg node1032_r;
    reg node1032_l;
    reg node1033;
    reg node1034;
    reg node1035_r;
    reg node1035_l;
    reg node1036;
    reg node1037;
    reg node1038_r;
    reg node1038_l;
    reg node1039_r;
    reg node1039_l;
    reg node1040_r;
    reg node1040_l;
    reg node1041_r;
    reg node1041_l;
    reg node1042_r;
    reg node1042_l;
    reg node1043;
    reg node1044;
    reg node1045_r;
    reg node1045_l;
    reg node1046;
    reg node1047;
    reg node1048_r;
    reg node1048_l;
    reg node1049_r;
    reg node1049_l;
    reg node1050;
    reg node1051;
    reg node1052_r;
    reg node1052_l;
    reg node1053;
    reg node1054;
    reg node1055_r;
    reg node1055_l;
    reg node1056_r;
    reg node1056_l;
    reg node1057;
    reg node1058;
    reg node1059;
    reg node1060_r;
    reg node1060_l;
    reg node1061_r;
    reg node1061_l;
    reg node1062_r;
    reg node1062_l;
    reg node1063_r;
    reg node1063_l;
    reg node1064;
    reg node1065;
    reg node1066_r;
    reg node1066_l;
    reg node1067;
    reg node1068;
    reg node1069_r;
    reg node1069_l;
    reg node1070_r;
    reg node1070_l;
    reg node1071;
    reg node1072;
    reg node1073_r;
    reg node1073_l;
    reg node1074;
    reg node1075;
    reg node1076_r;
    reg node1076_l;
    reg node1077_r;
    reg node1077_l;
    reg node1078_r;
    reg node1078_l;
    reg node1079;
    reg node1080;
    reg node1081_r;
    reg node1081_l;
    reg node1082;
    reg node1083;
    reg node1084_r;
    reg node1084_l;
    reg node1085_r;
    reg node1085_l;
    reg node1086;
    reg node1087;
    reg node1088_r;
    reg node1088_l;
    reg node1089;
    reg node1090;
    reg node1091_r;
    reg node1091_l;
    reg node1092_r;
    reg node1092_l;
    reg node1093_r;
    reg node1093_l;
    reg node1094_r;
    reg node1094_l;
    reg node1095_r;
    reg node1095_l;
    reg node1096_r;
    reg node1096_l;
    reg node1097_r;
    reg node1097_l;
    reg node1098;
    reg node1099;
    reg node1100_r;
    reg node1100_l;
    reg node1101;
    reg node1102;
    reg node1103_r;
    reg node1103_l;
    reg node1104_r;
    reg node1104_l;
    reg node1105;
    reg node1106;
    reg node1107;
    reg node1108_r;
    reg node1108_l;
    reg node1109_r;
    reg node1109_l;
    reg node1110_r;
    reg node1110_l;
    reg node1111;
    reg node1112;
    reg node1113_r;
    reg node1113_l;
    reg node1114;
    reg node1115;
    reg node1116_r;
    reg node1116_l;
    reg node1117_r;
    reg node1117_l;
    reg node1118;
    reg node1119;
    reg node1120_r;
    reg node1120_l;
    reg node1121;
    reg node1122;
    reg node1123_r;
    reg node1123_l;
    reg node1124_r;
    reg node1124_l;
    reg node1125_r;
    reg node1125_l;
    reg node1126_r;
    reg node1126_l;
    reg node1127;
    reg node1128;
    reg node1129_r;
    reg node1129_l;
    reg node1130;
    reg node1131;
    reg node1132_r;
    reg node1132_l;
    reg node1133_r;
    reg node1133_l;
    reg node1134;
    reg node1135;
    reg node1136;
    reg node1137_r;
    reg node1137_l;
    reg node1138_r;
    reg node1138_l;
    reg node1139_r;
    reg node1139_l;
    reg node1140;
    reg node1141;
    reg node1142_r;
    reg node1142_l;
    reg node1143;
    reg node1144;
    reg node1145_r;
    reg node1145_l;
    reg node1146_r;
    reg node1146_l;
    reg node1147;
    reg node1148;
    reg node1149_r;
    reg node1149_l;
    reg node1150;
    reg node1151;
    reg node1152_r;
    reg node1152_l;
    reg node1153_r;
    reg node1153_l;
    reg node1154_r;
    reg node1154_l;
    reg node1155_r;
    reg node1155_l;
    reg node1156_r;
    reg node1156_l;
    reg node1157;
    reg node1158;
    reg node1159_r;
    reg node1159_l;
    reg node1160;
    reg node1161;
    reg node1162_r;
    reg node1162_l;
    reg node1163_r;
    reg node1163_l;
    reg node1164;
    reg node1165;
    reg node1166_r;
    reg node1166_l;
    reg node1167;
    reg node1168;
    reg node1169_r;
    reg node1169_l;
    reg node1170_r;
    reg node1170_l;
    reg node1171_r;
    reg node1171_l;
    reg node1172;
    reg node1173;
    reg node1174_r;
    reg node1174_l;
    reg node1175;
    reg node1176;
    reg node1177_r;
    reg node1177_l;
    reg node1178;
    reg node1179_r;
    reg node1179_l;
    reg node1180;
    reg node1181;
    reg node1182_r;
    reg node1182_l;
    reg node1183_r;
    reg node1183_l;
    reg node1184_r;
    reg node1184_l;
    reg node1185_r;
    reg node1185_l;
    reg node1186;
    reg node1187;
    reg node1188_r;
    reg node1188_l;
    reg node1189;
    reg node1190;
    reg node1191_r;
    reg node1191_l;
    reg node1192_r;
    reg node1192_l;
    reg node1193;
    reg node1194;
    reg node1195_r;
    reg node1195_l;
    reg node1196;
    reg node1197;
    reg node1198_r;
    reg node1198_l;
    reg node1199_r;
    reg node1199_l;
    reg node1200_r;
    reg node1200_l;
    reg node1201;
    reg node1202;
    reg node1203_r;
    reg node1203_l;
    reg node1204;
    reg node1205;
    reg node1206_r;
    reg node1206_l;
    reg node1207_r;
    reg node1207_l;
    reg node1208;
    reg node1209;
    reg node1210_r;
    reg node1210_l;
    reg node1211;
    reg node1212;
    reg node1213_r;
    reg node1213_l;
    reg node1214_r;
    reg node1214_l;
    reg node1215_r;
    reg node1215_l;
    reg node1216_r;
    reg node1216_l;
    reg node1217_r;
    reg node1217_l;
    reg node1218_r;
    reg node1218_l;
    reg node1219;
    reg node1220;
    reg node1221_r;
    reg node1221_l;
    reg node1222;
    reg node1223;
    reg node1224_r;
    reg node1224_l;
    reg node1225_r;
    reg node1225_l;
    reg node1226;
    reg node1227;
    reg node1228;
    reg node1229_r;
    reg node1229_l;
    reg node1230_r;
    reg node1230_l;
    reg node1231_r;
    reg node1231_l;
    reg node1232;
    reg node1233;
    reg node1234_r;
    reg node1234_l;
    reg node1235;
    reg node1236;
    reg node1237_r;
    reg node1237_l;
    reg node1238_r;
    reg node1238_l;
    reg node1239;
    reg node1240;
    reg node1241;
    reg node1242_r;
    reg node1242_l;
    reg node1243_r;
    reg node1243_l;
    reg node1244_r;
    reg node1244_l;
    reg node1245_r;
    reg node1245_l;
    reg node1246;
    reg node1247;
    reg node1248_r;
    reg node1248_l;
    reg node1249;
    reg node1250;
    reg node1251_r;
    reg node1251_l;
    reg node1252_r;
    reg node1252_l;
    reg node1253;
    reg node1254;
    reg node1255_r;
    reg node1255_l;
    reg node1256;
    reg node1257;
    reg node1258_r;
    reg node1258_l;
    reg node1259_r;
    reg node1259_l;
    reg node1260_r;
    reg node1260_l;
    reg node1261;
    reg node1262;
    reg node1263;
    reg node1264_r;
    reg node1264_l;
    reg node1265_r;
    reg node1265_l;
    reg node1266;
    reg node1267;
    reg node1268;
    reg node1269_r;
    reg node1269_l;
    reg node1270_r;
    reg node1270_l;
    reg node1271_r;
    reg node1271_l;
    reg node1272_r;
    reg node1272_l;
    reg node1273;
    reg node1274_r;
    reg node1274_l;
    reg node1275;
    reg node1276;
    reg node1277_r;
    reg node1277_l;
    reg node1278;
    reg node1279_r;
    reg node1279_l;
    reg node1280;
    reg node1281;
    reg node1282_r;
    reg node1282_l;
    reg node1283_r;
    reg node1283_l;
    reg node1284;
    reg node1285;
    reg node1286_r;
    reg node1286_l;
    reg node1287;
    reg node1288_r;
    reg node1288_l;
    reg node1289;
    reg node1290;
    reg node1291_r;
    reg node1291_l;
    reg node1292_r;
    reg node1292_l;
    reg node1293_r;
    reg node1293_l;
    reg node1294_r;
    reg node1294_l;
    reg node1295;
    reg node1296;
    reg node1297_r;
    reg node1297_l;
    reg node1298;
    reg node1299;
    reg node1300_r;
    reg node1300_l;
    reg node1301;
    reg node1302;
    reg node1303_r;
    reg node1303_l;
    reg node1304_r;
    reg node1304_l;
    reg node1305;
    reg node1306;
    reg node1307_r;
    reg node1307_l;
    reg node1308_r;
    reg node1308_l;
    reg node1309;
    reg node1310;
    reg node1311;
    reg node1312_r;
    reg node1312_l;
    reg node1313_r;
    reg node1313_l;
    reg node1314_r;
    reg node1314_l;
    reg node1315_r;
    reg node1315_l;
    reg node1316_r;
    reg node1316_l;
    reg node1317_r;
    reg node1317_l;
    reg node1318_r;
    reg node1318_l;
    reg node1319_r;
    reg node1319_l;
    reg node1320;
    reg node1321;
    reg node1322;
    reg node1323_r;
    reg node1323_l;
    reg node1324_r;
    reg node1324_l;
    reg node1325;
    reg node1326;
    reg node1327;
    reg node1328_r;
    reg node1328_l;
    reg node1329_r;
    reg node1329_l;
    reg node1330_r;
    reg node1330_l;
    reg node1331;
    reg node1332;
    reg node1333;
    reg node1334_r;
    reg node1334_l;
    reg node1335_r;
    reg node1335_l;
    reg node1336;
    reg node1337;
    reg node1338;
    reg node1339_r;
    reg node1339_l;
    reg node1340_r;
    reg node1340_l;
    reg node1341_r;
    reg node1341_l;
    reg node1342_r;
    reg node1342_l;
    reg node1343;
    reg node1344;
    reg node1345_r;
    reg node1345_l;
    reg node1346;
    reg node1347;
    reg node1348_r;
    reg node1348_l;
    reg node1349_r;
    reg node1349_l;
    reg node1350;
    reg node1351;
    reg node1352_r;
    reg node1352_l;
    reg node1353;
    reg node1354;
    reg node1355_r;
    reg node1355_l;
    reg node1356_r;
    reg node1356_l;
    reg node1357_r;
    reg node1357_l;
    reg node1358;
    reg node1359;
    reg node1360;
    reg node1361_r;
    reg node1361_l;
    reg node1362;
    reg node1363_r;
    reg node1363_l;
    reg node1364;
    reg node1365;
    reg node1366_r;
    reg node1366_l;
    reg node1367_r;
    reg node1367_l;
    reg node1368_r;
    reg node1368_l;
    reg node1369_r;
    reg node1369_l;
    reg node1370_r;
    reg node1370_l;
    reg node1371;
    reg node1372;
    reg node1373;
    reg node1374_r;
    reg node1374_l;
    reg node1375_r;
    reg node1375_l;
    reg node1376;
    reg node1377;
    reg node1378_r;
    reg node1378_l;
    reg node1379;
    reg node1380;
    reg node1381_r;
    reg node1381_l;
    reg node1382_r;
    reg node1382_l;
    reg node1383_r;
    reg node1383_l;
    reg node1384;
    reg node1385;
    reg node1386_r;
    reg node1386_l;
    reg node1387;
    reg node1388;
    reg node1389_r;
    reg node1389_l;
    reg node1390_r;
    reg node1390_l;
    reg node1391;
    reg node1392;
    reg node1393_r;
    reg node1393_l;
    reg node1394;
    reg node1395;
    reg node1396_r;
    reg node1396_l;
    reg node1397_r;
    reg node1397_l;
    reg node1398_r;
    reg node1398_l;
    reg node1399_r;
    reg node1399_l;
    reg node1400;
    reg node1401;
    reg node1402;
    reg node1403_r;
    reg node1403_l;
    reg node1404;
    reg node1405;
    reg node1406_r;
    reg node1406_l;
    reg node1407_r;
    reg node1407_l;
    reg node1408_r;
    reg node1408_l;
    reg node1409;
    reg node1410;
    reg node1411_r;
    reg node1411_l;
    reg node1412;
    reg node1413;
    reg node1414_r;
    reg node1414_l;
    reg node1415;
    reg node1416;
    reg node1417_r;
    reg node1417_l;
    reg node1418_r;
    reg node1418_l;
    reg node1419_r;
    reg node1419_l;
    reg node1420_r;
    reg node1420_l;
    reg node1421_r;
    reg node1421_l;
    reg node1422_r;
    reg node1422_l;
    reg node1423;
    reg node1424;
    reg node1425_r;
    reg node1425_l;
    reg node1426;
    reg node1427;
    reg node1428_r;
    reg node1428_l;
    reg node1429_r;
    reg node1429_l;
    reg node1430;
    reg node1431;
    reg node1432_r;
    reg node1432_l;
    reg node1433;
    reg node1434;
    reg node1435_r;
    reg node1435_l;
    reg node1436_r;
    reg node1436_l;
    reg node1437_r;
    reg node1437_l;
    reg node1438;
    reg node1439;
    reg node1440_r;
    reg node1440_l;
    reg node1441;
    reg node1442;
    reg node1443_r;
    reg node1443_l;
    reg node1444_r;
    reg node1444_l;
    reg node1445;
    reg node1446;
    reg node1447;
    reg node1448_r;
    reg node1448_l;
    reg node1449_r;
    reg node1449_l;
    reg node1450_r;
    reg node1450_l;
    reg node1451_r;
    reg node1451_l;
    reg node1452;
    reg node1453;
    reg node1454_r;
    reg node1454_l;
    reg node1455;
    reg node1456;
    reg node1457_r;
    reg node1457_l;
    reg node1458;
    reg node1459_r;
    reg node1459_l;
    reg node1460;
    reg node1461;
    reg node1462_r;
    reg node1462_l;
    reg node1463_r;
    reg node1463_l;
    reg node1464_r;
    reg node1464_l;
    reg node1465;
    reg node1466;
    reg node1467;
    reg node1468_r;
    reg node1468_l;
    reg node1469;
    reg node1470_r;
    reg node1470_l;
    reg node1471;
    reg node1472;
    reg node1473_r;
    reg node1473_l;
    reg node1474_r;
    reg node1474_l;
    reg node1475_r;
    reg node1475_l;
    reg node1476_r;
    reg node1476_l;
    reg node1477_r;
    reg node1477_l;
    reg node1478;
    reg node1479;
    reg node1480;
    reg node1481_r;
    reg node1481_l;
    reg node1482;
    reg node1483;
    reg node1484_r;
    reg node1484_l;
    reg node1485_r;
    reg node1485_l;
    reg node1486;
    reg node1487;
    reg node1488_r;
    reg node1488_l;
    reg node1489_r;
    reg node1489_l;
    reg node1490;
    reg node1491;
    reg node1492_r;
    reg node1492_l;
    reg node1493;
    reg node1494;
    reg node1495_r;
    reg node1495_l;
    reg node1496_r;
    reg node1496_l;
    reg node1497_r;
    reg node1497_l;
    reg node1498_r;
    reg node1498_l;
    reg node1499;
    reg node1500;
    reg node1501_r;
    reg node1501_l;
    reg node1502;
    reg node1503;
    reg node1504_r;
    reg node1504_l;
    reg node1505_r;
    reg node1505_l;
    reg node1506;
    reg node1507;
    reg node1508_r;
    reg node1508_l;
    reg node1509;
    reg node1510;
    reg node1511_r;
    reg node1511_l;
    reg node1512_r;
    reg node1512_l;
    reg node1513_r;
    reg node1513_l;
    reg node1514;
    reg node1515;
    reg node1516_r;
    reg node1516_l;
    reg node1517;
    reg node1518;
    reg node1519_r;
    reg node1519_l;
    reg node1520_r;
    reg node1520_l;
    reg node1521;
    reg node1522;
    reg node1523;
    reg node1524_r;
    reg node1524_l;
    reg node1525_r;
    reg node1525_l;
    reg node1526_r;
    reg node1526_l;
    reg node1527_r;
    reg node1527_l;
    reg node1528_r;
    reg node1528_l;
    reg node1529_r;
    reg node1529_l;
    reg node1530_r;
    reg node1530_l;
    reg node1531;
    reg node1532;
    reg node1533_r;
    reg node1533_l;
    reg node1534;
    reg node1535;
    reg node1536_r;
    reg node1536_l;
    reg node1537_r;
    reg node1537_l;
    reg node1538;
    reg node1539;
    reg node1540_r;
    reg node1540_l;
    reg node1541;
    reg node1542;
    reg node1543_r;
    reg node1543_l;
    reg node1544_r;
    reg node1544_l;
    reg node1545_r;
    reg node1545_l;
    reg node1546;
    reg node1547;
    reg node1548_r;
    reg node1548_l;
    reg node1549;
    reg node1550;
    reg node1551_r;
    reg node1551_l;
    reg node1552_r;
    reg node1552_l;
    reg node1553;
    reg node1554;
    reg node1555_r;
    reg node1555_l;
    reg node1556;
    reg node1557;
    reg node1558_r;
    reg node1558_l;
    reg node1559_r;
    reg node1559_l;
    reg node1560_r;
    reg node1560_l;
    reg node1561_r;
    reg node1561_l;
    reg node1562;
    reg node1563;
    reg node1564_r;
    reg node1564_l;
    reg node1565;
    reg node1566;
    reg node1567_r;
    reg node1567_l;
    reg node1568_r;
    reg node1568_l;
    reg node1569;
    reg node1570;
    reg node1571_r;
    reg node1571_l;
    reg node1572;
    reg node1573;
    reg node1574_r;
    reg node1574_l;
    reg node1575_r;
    reg node1575_l;
    reg node1576_r;
    reg node1576_l;
    reg node1577;
    reg node1578;
    reg node1579_r;
    reg node1579_l;
    reg node1580;
    reg node1581;
    reg node1582_r;
    reg node1582_l;
    reg node1583_r;
    reg node1583_l;
    reg node1584;
    reg node1585;
    reg node1586_r;
    reg node1586_l;
    reg node1587;
    reg node1588;
    reg node1589_r;
    reg node1589_l;
    reg node1590_r;
    reg node1590_l;
    reg node1591_r;
    reg node1591_l;
    reg node1592_r;
    reg node1592_l;
    reg node1593_r;
    reg node1593_l;
    reg node1594;
    reg node1595;
    reg node1596_r;
    reg node1596_l;
    reg node1597;
    reg node1598;
    reg node1599_r;
    reg node1599_l;
    reg node1600_r;
    reg node1600_l;
    reg node1601;
    reg node1602;
    reg node1603_r;
    reg node1603_l;
    reg node1604;
    reg node1605;
    reg node1606_r;
    reg node1606_l;
    reg node1607;
    reg node1608_r;
    reg node1608_l;
    reg node1609;
    reg node1610_r;
    reg node1610_l;
    reg node1611;
    reg node1612;
    reg node1613_r;
    reg node1613_l;
    reg node1614_r;
    reg node1614_l;
    reg node1615_r;
    reg node1615_l;
    reg node1616_r;
    reg node1616_l;
    reg node1617;
    reg node1618;
    reg node1619_r;
    reg node1619_l;
    reg node1620;
    reg node1621;
    reg node1622;
    reg node1623_r;
    reg node1623_l;
    reg node1624;
    reg node1625_r;
    reg node1625_l;
    reg node1626;
    reg node1627_r;
    reg node1627_l;
    reg node1628;
    reg node1629;
    reg node1630_r;
    reg node1630_l;
    reg node1631_r;
    reg node1631_l;
    reg node1632_r;
    reg node1632_l;
    reg node1633_r;
    reg node1633_l;
    reg node1634_r;
    reg node1634_l;
    reg node1635_r;
    reg node1635_l;
    reg node1636;
    reg node1637;
    reg node1638_r;
    reg node1638_l;
    reg node1639;
    reg node1640;
    reg node1641_r;
    reg node1641_l;
    reg node1642_r;
    reg node1642_l;
    reg node1643;
    reg node1644;
    reg node1645;
    reg node1646_r;
    reg node1646_l;
    reg node1647_r;
    reg node1647_l;
    reg node1648_r;
    reg node1648_l;
    reg node1649;
    reg node1650;
    reg node1651_r;
    reg node1651_l;
    reg node1652;
    reg node1653;
    reg node1654_r;
    reg node1654_l;
    reg node1655_r;
    reg node1655_l;
    reg node1656;
    reg node1657;
    reg node1658_r;
    reg node1658_l;
    reg node1659;
    reg node1660;
    reg node1661_r;
    reg node1661_l;
    reg node1662_r;
    reg node1662_l;
    reg node1663_r;
    reg node1663_l;
    reg node1664_r;
    reg node1664_l;
    reg node1665;
    reg node1666;
    reg node1667_r;
    reg node1667_l;
    reg node1668;
    reg node1669;
    reg node1670;
    reg node1671_r;
    reg node1671_l;
    reg node1672_r;
    reg node1672_l;
    reg node1673_r;
    reg node1673_l;
    reg node1674;
    reg node1675;
    reg node1676;
    reg node1677_r;
    reg node1677_l;
    reg node1678_r;
    reg node1678_l;
    reg node1679;
    reg node1680;
    reg node1681_r;
    reg node1681_l;
    reg node1682;
    reg node1683;
    reg node1684_r;
    reg node1684_l;
    reg node1685_r;
    reg node1685_l;
    reg node1686_r;
    reg node1686_l;
    reg node1687_r;
    reg node1687_l;
    reg node1688_r;
    reg node1688_l;
    reg node1689;
    reg node1690;
    reg node1691_r;
    reg node1691_l;
    reg node1692;
    reg node1693;
    reg node1694_r;
    reg node1694_l;
    reg node1695_r;
    reg node1695_l;
    reg node1696;
    reg node1697;
    reg node1698_r;
    reg node1698_l;
    reg node1699;
    reg node1700;
    reg node1701_r;
    reg node1701_l;
    reg node1702_r;
    reg node1702_l;
    reg node1703_r;
    reg node1703_l;
    reg node1704;
    reg node1705;
    reg node1706_r;
    reg node1706_l;
    reg node1707;
    reg node1708;
    reg node1709_r;
    reg node1709_l;
    reg node1710_r;
    reg node1710_l;
    reg node1711;
    reg node1712;
    reg node1713_r;
    reg node1713_l;
    reg node1714;
    reg node1715;
    reg node1716_r;
    reg node1716_l;
    reg node1717_r;
    reg node1717_l;
    reg node1718;
    reg node1719;
    reg node1720_r;
    reg node1720_l;
    reg node1721;
    reg node1722_r;
    reg node1722_l;
    reg node1723;
    reg node1724;
    reg result0;
    reg result1;
    reg result2;
    reg result3;
    reg result4;
    reg result5;
    reg result6;
    reg result7;
    reg result8;
    reg result9;

    begin
      node0_r = pixel[541];
      node0_l = ~pixel[541];
      node1_r = node0_l & pixel[437];
      node1_l = node0_l & ~pixel[437];
      node2_r = node1_l & pixel[454];
      node2_l = node1_l & ~pixel[454];
      node3_r = node2_l & pixel[347];
      node3_l = node2_l & ~pixel[347];
      node4_r = node3_l & pixel[262];
      node4_l = node3_l & ~pixel[262];
      node5_r = node4_l & pixel[578];
      node5_l = node4_l & ~pixel[578];
      node6_r = node5_l & pixel[458];
      node6_l = node5_l & ~pixel[458];
      node7_r = node6_l & pixel[233];
      node7_l = node6_l & ~pixel[233];
      node8_r = node7_l & pixel[327];
      node8_l = node7_l & ~pixel[327];
      node9_r = node8_l & pixel[175];
      node9_l = node8_l & ~pixel[175];
      node10 = node9_l;
      node11 = node9_r;
      node12_r = node8_r & pixel[292];
      node12_l = node8_r & ~pixel[292];
      node13 = node12_l;
      node14 = node12_r;
      node15_r = node7_r & pixel[636];
      node15_l = node7_r & ~pixel[636];
      node16_r = node15_l & pixel[124];
      node16_l = node15_l & ~pixel[124];
      node17 = node16_l;
      node18 = node16_r;
      node19_r = node15_r & pixel[525];
      node19_l = node15_r & ~pixel[525];
      node20 = node19_l;
      node21 = node19_r;
      node22_r = node6_r & pixel[180];
      node22_l = node6_r & ~pixel[180];
      node23_r = node22_l & pixel[219];
      node23_l = node22_l & ~pixel[219];
      node24_r = node23_l & pixel[567];
      node24_l = node23_l & ~pixel[567];
      node25 = node24_l;
      node26 = node24_r;
      node27_r = node23_r & pixel[345];
      node27_l = node23_r & ~pixel[345];
      node28 = node27_l;
      node29 = node27_r;
      node30_r = node22_r & pixel[430];
      node30_l = node22_r & ~pixel[430];
      node31_r = node30_l & pixel[600];
      node31_l = node30_l & ~pixel[600];
      node32 = node31_l;
      node33 = node31_r;
      node34_r = node30_r & pixel[539];
      node34_l = node30_r & ~pixel[539];
      node35 = node34_l;
      node36 = node34_r;
      node37_r = node5_r & pixel[543];
      node37_l = node5_r & ~pixel[543];
      node38_r = node37_l & pixel[320];
      node38_l = node37_l & ~pixel[320];
      node39_r = node38_l & pixel[658];
      node39_l = node38_l & ~pixel[658];
      node40_r = node39_l & pixel[512];
      node40_l = node39_l & ~pixel[512];
      node41 = node40_l;
      node42 = node40_r;
      node43_r = node39_r & pixel[582];
      node43_l = node39_r & ~pixel[582];
      node44 = node43_l;
      node45 = node43_r;
      node46_r = node38_r & pixel[325];
      node46_l = node38_r & ~pixel[325];
      node47_r = node46_l & pixel[215];
      node47_l = node46_l & ~pixel[215];
      node48 = node47_l;
      node49 = node47_r;
      node50_r = node46_r & pixel[435];
      node50_l = node46_r & ~pixel[435];
      node51 = node50_l;
      node52 = node50_r;
      node53_r = node37_r & pixel[345];
      node53_l = node37_r & ~pixel[345];
      node54_r = node53_l & pixel[456];
      node54_l = node53_l & ~pixel[456];
      node55_r = node54_l & pixel[348];
      node55_l = node54_l & ~pixel[348];
      node56 = node55_l;
      node57 = node55_r;
      node58 = node54_r;
      node59_r = node53_r & pixel[153];
      node59_l = node53_r & ~pixel[153];
      node60 = node59_l;
      node61_r = node59_r & pixel[185];
      node61_l = node59_r & ~pixel[185];
      node62 = node61_l;
      node63 = node61_r;
      node64_r = node4_r & pixel[429];
      node64_l = node4_r & ~pixel[429];
      node65_r = node64_l & pixel[183];
      node65_l = node64_l & ~pixel[183];
      node66_r = node65_l & pixel[555];
      node66_l = node65_l & ~pixel[555];
      node67_r = node66_l & pixel[402];
      node67_l = node66_l & ~pixel[402];
      node68_r = node67_l & pixel[604];
      node68_l = node67_l & ~pixel[604];
      node69 = node68_l;
      node70 = node68_r;
      node71_r = node67_r & pixel[523];
      node71_l = node67_r & ~pixel[523];
      node72 = node71_l;
      node73 = node71_r;
      node74_r = node66_r & pixel[433];
      node74_l = node66_r & ~pixel[433];
      node75 = node74_l;
      node76_r = node74_r & pixel[546];
      node76_l = node74_r & ~pixel[546];
      node77 = node76_l;
      node78 = node76_r;
      node79_r = node65_r & pixel[681];
      node79_l = node65_r & ~pixel[681];
      node80_r = node79_l & pixel[404];
      node80_l = node79_l & ~pixel[404];
      node81_r = node80_l & pixel[154];
      node81_l = node80_l & ~pixel[154];
      node82 = node81_l;
      node83 = node81_r;
      node84_r = node80_r & pixel[472];
      node84_l = node80_r & ~pixel[472];
      node85 = node84_l;
      node86 = node84_r;
      node87_r = node79_r & pixel[545];
      node87_l = node79_r & ~pixel[545];
      node88_r = node87_l & pixel[379];
      node88_l = node87_l & ~pixel[379];
      node89 = node88_l;
      node90 = node88_r;
      node91_r = node87_r & pixel[544];
      node91_l = node87_r & ~pixel[544];
      node92 = node91_l;
      node93 = node91_r;
      node94_r = node64_r & pixel[238];
      node94_l = node64_r & ~pixel[238];
      node95_r = node94_l & pixel[572];
      node95_l = node94_l & ~pixel[572];
      node96_r = node95_l & pixel[321];
      node96_l = node95_l & ~pixel[321];
      node97_r = node96_l & pixel[298];
      node97_l = node96_l & ~pixel[298];
      node98 = node97_l;
      node99 = node97_r;
      node100_r = node96_r & pixel[718];
      node100_l = node96_r & ~pixel[718];
      node101 = node100_l;
      node102 = node100_r;
      node103_r = node95_r & pixel[657];
      node103_l = node95_r & ~pixel[657];
      node104_r = node103_l & pixel[398];
      node104_l = node103_l & ~pixel[398];
      node105 = node104_l;
      node106 = node104_r;
      node107_r = node103_r & pixel[380];
      node107_l = node103_r & ~pixel[380];
      node108 = node107_l;
      node109 = node107_r;
      node110_r = node94_r & pixel[324];
      node110_l = node94_r & ~pixel[324];
      node111_r = node110_l & pixel[317];
      node111_l = node110_l & ~pixel[317];
      node112_r = node111_l & pixel[438];
      node112_l = node111_l & ~pixel[438];
      node113 = node112_l;
      node114 = node112_r;
      node115_r = node111_r & pixel[325];
      node115_l = node111_r & ~pixel[325];
      node116 = node115_l;
      node117 = node115_r;
      node118_r = node110_r & pixel[155];
      node118_l = node110_r & ~pixel[155];
      node119_r = node118_l & pixel[289];
      node119_l = node118_l & ~pixel[289];
      node120 = node119_l;
      node121 = node119_r;
      node122_r = node118_r & pixel[441];
      node122_l = node118_r & ~pixel[441];
      node123 = node122_l;
      node124 = node122_r;
      node125_r = node3_r & pixel[220];
      node125_l = node3_r & ~pixel[220];
      node126_r = node125_l & pixel[435];
      node126_l = node125_l & ~pixel[435];
      node127_r = node126_l & pixel[290];
      node127_l = node126_l & ~pixel[290];
      node128_r = node127_l & pixel[496];
      node128_l = node127_l & ~pixel[496];
      node129_r = node128_l & pixel[468];
      node129_l = node128_l & ~pixel[468];
      node130_r = node129_l & pixel[542];
      node130_l = node129_l & ~pixel[542];
      node131 = node130_l;
      node132 = node130_r;
      node133_r = node129_r & pixel[328];
      node133_l = node129_r & ~pixel[328];
      node134 = node133_l;
      node135 = node133_r;
      node136_r = node128_r & pixel[154];
      node136_l = node128_r & ~pixel[154];
      node137_r = node136_l & pixel[351];
      node137_l = node136_l & ~pixel[351];
      node138 = node137_l;
      node139 = node137_r;
      node140_r = node136_r & pixel[289];
      node140_l = node136_r & ~pixel[289];
      node141 = node140_l;
      node142 = node140_r;
      node143_r = node127_r & pixel[403];
      node143_l = node127_r & ~pixel[403];
      node144_r = node143_l & pixel[284];
      node144_l = node143_l & ~pixel[284];
      node145_r = node144_l & pixel[428];
      node145_l = node144_l & ~pixel[428];
      node146 = node145_l;
      node147 = node145_r;
      node148_r = node144_r & pixel[155];
      node148_l = node144_r & ~pixel[155];
      node149 = node148_l;
      node150 = node148_r;
      node151_r = node143_r & pixel[657];
      node151_l = node143_r & ~pixel[657];
      node152_r = node151_l & pixel[606];
      node152_l = node151_l & ~pixel[606];
      node153 = node152_l;
      node154 = node152_r;
      node155_r = node151_r & pixel[382];
      node155_l = node151_r & ~pixel[382];
      node156 = node155_l;
      node157 = node155_r;
      node158_r = node126_r & pixel[521];
      node158_l = node126_r & ~pixel[521];
      node159_r = node158_l & pixel[154];
      node159_l = node158_l & ~pixel[154];
      node160_r = node159_l & pixel[211];
      node160_l = node159_l & ~pixel[211];
      node161_r = node160_l & pixel[379];
      node161_l = node160_l & ~pixel[379];
      node162 = node161_l;
      node163 = node161_r;
      node164_r = node160_r & pixel[301];
      node164_l = node160_r & ~pixel[301];
      node165 = node164_l;
      node166 = node164_r;
      node167_r = node159_r & pixel[270];
      node167_l = node159_r & ~pixel[270];
      node168_r = node167_l & pixel[266];
      node168_l = node167_l & ~pixel[266];
      node169 = node168_l;
      node170 = node168_r;
      node171_r = node167_r & pixel[441];
      node171_l = node167_r & ~pixel[441];
      node172 = node171_l;
      node173 = node171_r;
      node174_r = node158_r & pixel[381];
      node174_l = node158_r & ~pixel[381];
      node175_r = node174_l & pixel[544];
      node175_l = node174_l & ~pixel[544];
      node176_r = node175_l & pixel[318];
      node176_l = node175_l & ~pixel[318];
      node177 = node176_l;
      node178 = node176_r;
      node179_r = node175_r & pixel[127];
      node179_l = node175_r & ~pixel[127];
      node180 = node179_l;
      node181 = node179_r;
      node182_r = node174_r & pixel[383];
      node182_l = node174_r & ~pixel[383];
      node183_r = node182_l & pixel[605];
      node183_l = node182_l & ~pixel[605];
      node184 = node183_l;
      node185 = node183_r;
      node186_r = node182_r & pixel[329];
      node186_l = node182_r & ~pixel[329];
      node187 = node186_l;
      node188 = node186_r;
      node189_r = node125_r & pixel[511];
      node189_l = node125_r & ~pixel[511];
      node190_r = node189_l & pixel[353];
      node190_l = node189_l & ~pixel[353];
      node191 = node190_l;
      node192_r = node190_r & pixel[566];
      node192_l = node190_r & ~pixel[566];
      node193_r = node192_l & pixel[489];
      node193_l = node192_l & ~pixel[489];
      node194 = node193_l;
      node195_r = node193_r & pixel[288];
      node195_l = node193_r & ~pixel[288];
      node196 = node195_l;
      node197 = node195_r;
      node198 = node192_r;
      node199_r = node189_r & pixel[650];
      node199_l = node189_r & ~pixel[650];
      node200_r = node199_l & pixel[355];
      node200_l = node199_l & ~pixel[355];
      node201_r = node200_l & pixel[185];
      node201_l = node200_l & ~pixel[185];
      node202 = node201_l;
      node203_r = node201_r & pixel[326];
      node203_l = node201_r & ~pixel[326];
      node204 = node203_l;
      node205 = node203_r;
      node206_r = node200_r & pixel[430];
      node206_l = node200_r & ~pixel[430];
      node207 = node206_l;
      node208 = node206_r;
      node209_r = node199_r & pixel[467];
      node209_l = node199_r & ~pixel[467];
      node210_r = node209_l & pixel[353];
      node210_l = node209_l & ~pixel[353];
      node211_r = node210_l & pixel[577];
      node211_l = node210_l & ~pixel[577];
      node212 = node211_l;
      node213 = node211_r;
      node214_r = node210_r & pixel[579];
      node214_l = node210_r & ~pixel[579];
      node215 = node214_l;
      node216 = node214_r;
      node217 = node209_r;
      node218_r = node2_r & pixel[358];
      node218_l = node2_r & ~pixel[358];
      node219_r = node218_l & pixel[623];
      node219_l = node218_l & ~pixel[623];
      node220_r = node219_l & pixel[658];
      node220_l = node219_l & ~pixel[658];
      node221_r = node220_l & pixel[458];
      node221_l = node220_l & ~pixel[458];
      node222_r = node221_l & pixel[662];
      node222_l = node221_l & ~pixel[662];
      node223_r = node222_l & pixel[322];
      node223_l = node222_l & ~pixel[322];
      node224_r = node223_l & pixel[569];
      node224_l = node223_l & ~pixel[569];
      node225 = node224_l;
      node226 = node224_r;
      node227_r = node223_r & pixel[428];
      node227_l = node223_r & ~pixel[428];
      node228 = node227_l;
      node229 = node227_r;
      node230_r = node222_r & pixel[374];
      node230_l = node222_r & ~pixel[374];
      node231_r = node230_l & pixel[403];
      node231_l = node230_l & ~pixel[403];
      node232 = node231_l;
      node233 = node231_r;
      node234_r = node230_r & pixel[481];
      node234_l = node230_r & ~pixel[481];
      node235 = node234_l;
      node236 = node234_r;
      node237_r = node221_r & pixel[287];
      node237_l = node221_r & ~pixel[287];
      node238_r = node237_l & pixel[459];
      node238_l = node237_l & ~pixel[459];
      node239_r = node238_l & pixel[398];
      node239_l = node238_l & ~pixel[398];
      node240 = node239_l;
      node241 = node239_r;
      node242_r = node238_r & pixel[571];
      node242_l = node238_r & ~pixel[571];
      node243 = node242_l;
      node244 = node242_r;
      node245_r = node237_r & pixel[720];
      node245_l = node237_r & ~pixel[720];
      node246_r = node245_l & pixel[263];
      node246_l = node245_l & ~pixel[263];
      node247 = node246_l;
      node248 = node246_r;
      node249 = node245_r;
      node250_r = node220_r & pixel[540];
      node250_l = node220_r & ~pixel[540];
      node251_r = node250_l & pixel[268];
      node251_l = node250_l & ~pixel[268];
      node252_r = node251_l & pixel[302];
      node252_l = node251_l & ~pixel[302];
      node253_r = node252_l & pixel[495];
      node253_l = node252_l & ~pixel[495];
      node254 = node253_l;
      node255 = node253_r;
      node256 = node252_r;
      node257_r = node251_r & pixel[245];
      node257_l = node251_r & ~pixel[245];
      node258_r = node257_l & pixel[399];
      node258_l = node257_l & ~pixel[399];
      node259 = node258_l;
      node260 = node258_r;
      node261 = node257_r;
      node262_r = node250_r & pixel[380];
      node262_l = node250_r & ~pixel[380];
      node263 = node262_l;
      node264_r = node262_r & pixel[406];
      node264_l = node262_r & ~pixel[406];
      node265 = node264_l;
      node266 = node264_r;
      node267_r = node219_r & pixel[354];
      node267_l = node219_r & ~pixel[354];
      node268_r = node267_l & pixel[376];
      node268_l = node267_l & ~pixel[376];
      node269_r = node268_l & pixel[383];
      node269_l = node268_l & ~pixel[383];
      node270 = node269_l;
      node271_r = node269_r & pixel[400];
      node271_l = node269_r & ~pixel[400];
      node272_r = node271_l & pixel[153];
      node272_l = node271_l & ~pixel[153];
      node273 = node272_l;
      node274 = node272_r;
      node275_r = node271_r & pixel[655];
      node275_l = node271_r & ~pixel[655];
      node276 = node275_l;
      node277 = node275_r;
      node278_r = node268_r & pixel[429];
      node278_l = node268_r & ~pixel[429];
      node279_r = node278_l & pixel[236];
      node279_l = node278_l & ~pixel[236];
      node280 = node279_l;
      node281_r = node279_r & pixel[527];
      node281_l = node279_r & ~pixel[527];
      node282 = node281_l;
      node283 = node281_r;
      node284_r = node278_r & pixel[511];
      node284_l = node278_r & ~pixel[511];
      node285_r = node284_l & pixel[413];
      node285_l = node284_l & ~pixel[413];
      node286 = node285_l;
      node287 = node285_r;
      node288 = node284_r;
      node289_r = node267_r & pixel[151];
      node289_l = node267_r & ~pixel[151];
      node290_r = node289_l & pixel[344];
      node290_l = node289_l & ~pixel[344];
      node291_r = node290_l & pixel[431];
      node291_l = node290_l & ~pixel[431];
      node292_r = node291_l & pixel[563];
      node292_l = node291_l & ~pixel[563];
      node293 = node292_l;
      node294 = node292_r;
      node295_r = node291_r & pixel[407];
      node295_l = node291_r & ~pixel[407];
      node296 = node295_l;
      node297 = node295_r;
      node298_r = node290_r & pixel[327];
      node298_l = node290_r & ~pixel[327];
      node299 = node298_l;
      node300_r = node298_r & pixel[381];
      node300_l = node298_r & ~pixel[381];
      node301 = node300_l;
      node302 = node300_r;
      node303_r = node289_r & pixel[691];
      node303_l = node289_r & ~pixel[691];
      node304_r = node303_l & pixel[205];
      node304_l = node303_l & ~pixel[205];
      node305 = node304_l;
      node306_r = node304_r & pixel[238];
      node306_l = node304_r & ~pixel[238];
      node307 = node306_l;
      node308 = node306_r;
      node309_r = node303_r & pixel[651];
      node309_l = node303_r & ~pixel[651];
      node310 = node309_l;
      node311 = node309_r;
      node312_r = node218_r & pixel[461];
      node312_l = node218_r & ~pixel[461];
      node313_r = node312_l & pixel[187];
      node313_l = node312_l & ~pixel[187];
      node314_r = node313_l & pixel[627];
      node314_l = node313_l & ~pixel[627];
      node315_r = node314_l & pixel[486];
      node315_l = node314_l & ~pixel[486];
      node316_r = node315_l & pixel[595];
      node316_l = node315_l & ~pixel[595];
      node317_r = node316_l & pixel[377];
      node317_l = node316_l & ~pixel[377];
      node318 = node317_l;
      node319 = node317_r;
      node320 = node316_r;
      node321_r = node315_r & pixel[718];
      node321_l = node315_r & ~pixel[718];
      node322_r = node321_l & pixel[235];
      node322_l = node321_l & ~pixel[235];
      node323 = node322_l;
      node324 = node322_r;
      node325 = node321_r;
      node326_r = node314_r & pixel[352];
      node326_l = node314_r & ~pixel[352];
      node327_r = node326_l & pixel[509];
      node327_l = node326_l & ~pixel[509];
      node328_r = node327_l & pixel[482];
      node328_l = node327_l & ~pixel[482];
      node329 = node328_l;
      node330 = node328_r;
      node331 = node327_r;
      node332_r = node326_r & pixel[377];
      node332_l = node326_r & ~pixel[377];
      node333 = node332_l;
      node334_r = node332_r & pixel[270];
      node334_l = node332_r & ~pixel[270];
      node335 = node334_l;
      node336 = node334_r;
      node337_r = node313_r & pixel[380];
      node337_l = node313_r & ~pixel[380];
      node338_r = node337_l & pixel[352];
      node338_l = node337_l & ~pixel[352];
      node339_r = node338_l & pixel[407];
      node339_l = node338_l & ~pixel[407];
      node340_r = node339_l & pixel[174];
      node340_l = node339_l & ~pixel[174];
      node341 = node340_l;
      node342 = node340_r;
      node343_r = node339_r & pixel[290];
      node343_l = node339_r & ~pixel[290];
      node344 = node343_l;
      node345 = node343_r;
      node346_r = node338_r & pixel[214];
      node346_l = node338_r & ~pixel[214];
      node347 = node346_l;
      node348_r = node346_r & pixel[359];
      node348_l = node346_r & ~pixel[359];
      node349 = node348_l;
      node350 = node348_r;
      node351_r = node337_r & pixel[354];
      node351_l = node337_r & ~pixel[354];
      node352 = node351_l;
      node353_r = node351_r & pixel[547];
      node353_l = node351_r & ~pixel[547];
      node354_r = node353_l & pixel[404];
      node354_l = node353_l & ~pixel[404];
      node355 = node354_l;
      node356 = node354_r;
      node357_r = node353_r & pixel[235];
      node357_l = node353_r & ~pixel[235];
      node358 = node357_l;
      node359 = node357_r;
      node360_r = node312_r & pixel[345];
      node360_l = node312_r & ~pixel[345];
      node361_r = node360_l & pixel[353];
      node361_l = node360_l & ~pixel[353];
      node362_r = node361_l & pixel[567];
      node362_l = node361_l & ~pixel[567];
      node363_r = node362_l & pixel[286];
      node363_l = node362_l & ~pixel[286];
      node364_r = node363_l & pixel[217];
      node364_l = node363_l & ~pixel[217];
      node365 = node364_l;
      node366 = node364_r;
      node367 = node363_r;
      node368_r = node362_r & pixel[412];
      node368_l = node362_r & ~pixel[412];
      node369 = node368_l;
      node370 = node368_r;
      node371_r = node361_r & pixel[331];
      node371_l = node361_r & ~pixel[331];
      node372_r = node371_l & pixel[236];
      node372_l = node371_l & ~pixel[236];
      node373 = node372_l;
      node374 = node372_r;
      node375_r = node371_r & pixel[623];
      node375_l = node371_r & ~pixel[623];
      node376_r = node375_l & pixel[240];
      node376_l = node375_l & ~pixel[240];
      node377 = node376_l;
      node378 = node376_r;
      node379_r = node375_r & pixel[233];
      node379_l = node375_r & ~pixel[233];
      node380 = node379_l;
      node381 = node379_r;
      node382_r = node360_r & pixel[214];
      node382_l = node360_r & ~pixel[214];
      node383_r = node382_l & pixel[150];
      node383_l = node382_l & ~pixel[150];
      node384 = node383_l;
      node385_r = node383_r & pixel[128];
      node385_l = node383_r & ~pixel[128];
      node386 = node385_l;
      node387 = node385_r;
      node388_r = node382_r & pixel[713];
      node388_l = node382_r & ~pixel[713];
      node389_r = node388_l & pixel[369];
      node389_l = node388_l & ~pixel[369];
      node390 = node389_l;
      node391_r = node389_r & pixel[157];
      node391_l = node389_r & ~pixel[157];
      node392 = node391_l;
      node393 = node391_r;
      node394_r = node388_r & pixel[524];
      node394_l = node388_r & ~pixel[524];
      node395 = node394_l;
      node396 = node394_r;
      node397_r = node1_r & pixel[376];
      node397_l = node1_r & ~pixel[376];
      node398_r = node397_l & pixel[212];
      node398_l = node397_l & ~pixel[212];
      node399_r = node398_l & pixel[459];
      node399_l = node398_l & ~pixel[459];
      node400_r = node399_l & pixel[128];
      node400_l = node399_l & ~pixel[128];
      node401_r = node400_l & pixel[429];
      node401_l = node400_l & ~pixel[429];
      node402_r = node401_l & pixel[483];
      node402_l = node401_l & ~pixel[483];
      node403_r = node402_l & pixel[377];
      node403_l = node402_l & ~pixel[377];
      node404_r = node403_l & pixel[430];
      node404_l = node403_l & ~pixel[430];
      node405 = node404_l;
      node406 = node404_r;
      node407_r = node403_r & pixel[545];
      node407_l = node403_r & ~pixel[545];
      node408 = node407_l;
      node409 = node407_r;
      node410_r = node402_r & pixel[487];
      node410_l = node402_r & ~pixel[487];
      node411_r = node410_l & pixel[266];
      node411_l = node410_l & ~pixel[266];
      node412 = node411_l;
      node413 = node411_r;
      node414_r = node410_r & pixel[575];
      node414_l = node410_r & ~pixel[575];
      node415 = node414_l;
      node416 = node414_r;
      node417_r = node401_r & pixel[525];
      node417_l = node401_r & ~pixel[525];
      node418_r = node417_l & pixel[293];
      node418_l = node417_l & ~pixel[293];
      node419_r = node418_l & pixel[210];
      node419_l = node418_l & ~pixel[210];
      node420 = node419_l;
      node421 = node419_r;
      node422_r = node418_r & pixel[431];
      node422_l = node418_r & ~pixel[431];
      node423 = node422_l;
      node424 = node422_r;
      node425_r = node417_r & pixel[457];
      node425_l = node417_r & ~pixel[457];
      node426_r = node425_l & pixel[271];
      node426_l = node425_l & ~pixel[271];
      node427 = node426_l;
      node428 = node426_r;
      node429_r = node425_r & pixel[451];
      node429_l = node425_r & ~pixel[451];
      node430 = node429_l;
      node431 = node429_r;
      node432_r = node400_r & pixel[518];
      node432_l = node400_r & ~pixel[518];
      node433_r = node432_l & pixel[566];
      node433_l = node432_l & ~pixel[566];
      node434_r = node433_l & pixel[297];
      node434_l = node433_l & ~pixel[297];
      node435_r = node434_l & pixel[266];
      node435_l = node434_l & ~pixel[266];
      node436 = node435_l;
      node437 = node435_r;
      node438_r = node434_r & pixel[210];
      node438_l = node434_r & ~pixel[210];
      node439 = node438_l;
      node440 = node438_r;
      node441_r = node433_r & pixel[455];
      node441_l = node433_r & ~pixel[455];
      node442_r = node441_l & pixel[299];
      node442_l = node441_l & ~pixel[299];
      node443 = node442_l;
      node444 = node442_r;
      node445_r = node441_r & pixel[149];
      node445_l = node441_r & ~pixel[149];
      node446 = node445_l;
      node447 = node445_r;
      node448_r = node432_r & pixel[344];
      node448_l = node432_r & ~pixel[344];
      node449_r = node448_l & pixel[244];
      node449_l = node448_l & ~pixel[244];
      node450_r = node449_l & pixel[607];
      node450_l = node449_l & ~pixel[607];
      node451 = node450_l;
      node452 = node450_r;
      node453 = node449_r;
      node454_r = node448_r & pixel[347];
      node454_l = node448_r & ~pixel[347];
      node455 = node454_l;
      node456 = node454_r;
      node457_r = node399_r & pixel[239];
      node457_l = node399_r & ~pixel[239];
      node458_r = node457_l & pixel[128];
      node458_l = node457_l & ~pixel[128];
      node459_r = node458_l & pixel[322];
      node459_l = node458_l & ~pixel[322];
      node460_r = node459_l & pixel[460];
      node460_l = node459_l & ~pixel[460];
      node461_r = node460_l & pixel[426];
      node461_l = node460_l & ~pixel[426];
      node462 = node461_l;
      node463 = node461_r;
      node464_r = node460_r & pixel[498];
      node464_l = node460_r & ~pixel[498];
      node465 = node464_l;
      node466 = node464_r;
      node467_r = node459_r & pixel[161];
      node467_l = node459_r & ~pixel[161];
      node468_r = node467_l & pixel[552];
      node468_l = node467_l & ~pixel[552];
      node469 = node468_l;
      node470 = node468_r;
      node471_r = node467_r & pixel[629];
      node471_l = node467_r & ~pixel[629];
      node472 = node471_l;
      node473 = node471_r;
      node474_r = node458_r & pixel[539];
      node474_l = node458_r & ~pixel[539];
      node475_r = node474_l & pixel[508];
      node475_l = node474_l & ~pixel[508];
      node476_r = node475_l & pixel[657];
      node476_l = node475_l & ~pixel[657];
      node477 = node476_l;
      node478 = node476_r;
      node479_r = node475_r & pixel[656];
      node479_l = node475_r & ~pixel[656];
      node480 = node479_l;
      node481 = node479_r;
      node482_r = node474_r & pixel[374];
      node482_l = node474_r & ~pixel[374];
      node483_r = node482_l & pixel[323];
      node483_l = node482_l & ~pixel[323];
      node484 = node483_l;
      node485 = node483_r;
      node486_r = node482_r & pixel[465];
      node486_l = node482_r & ~pixel[465];
      node487 = node486_l;
      node488 = node486_r;
      node489_r = node457_r & pixel[347];
      node489_l = node457_r & ~pixel[347];
      node490_r = node489_l & pixel[602];
      node490_l = node489_l & ~pixel[602];
      node491_r = node490_l & pixel[409];
      node491_l = node490_l & ~pixel[409];
      node492_r = node491_l & pixel[151];
      node492_l = node491_l & ~pixel[151];
      node493 = node492_l;
      node494 = node492_r;
      node495_r = node491_r & pixel[208];
      node495_l = node491_r & ~pixel[208];
      node496 = node495_l;
      node497 = node495_r;
      node498_r = node490_r & pixel[258];
      node498_l = node490_r & ~pixel[258];
      node499_r = node498_l & pixel[203];
      node499_l = node498_l & ~pixel[203];
      node500 = node499_l;
      node501 = node499_r;
      node502_r = node498_r & pixel[397];
      node502_l = node498_r & ~pixel[397];
      node503 = node502_l;
      node504 = node502_r;
      node505_r = node489_r & pixel[261];
      node505_l = node489_r & ~pixel[261];
      node506_r = node505_l & pixel[210];
      node506_l = node505_l & ~pixel[210];
      node507_r = node506_l & pixel[595];
      node507_l = node506_l & ~pixel[595];
      node508 = node507_l;
      node509 = node507_r;
      node510_r = node506_r & pixel[130];
      node510_l = node506_r & ~pixel[130];
      node511 = node510_l;
      node512 = node510_r;
      node513_r = node505_r & pixel[256];
      node513_l = node505_r & ~pixel[256];
      node514_r = node513_l & pixel[400];
      node514_l = node513_l & ~pixel[400];
      node515 = node514_l;
      node516 = node514_r;
      node517 = node513_r;
      node518_r = node398_r & pixel[457];
      node518_l = node398_r & ~pixel[457];
      node519_r = node518_l & pixel[154];
      node519_l = node518_l & ~pixel[154];
      node520_r = node519_l & pixel[429];
      node520_l = node519_l & ~pixel[429];
      node521_r = node520_l & pixel[405];
      node521_l = node520_l & ~pixel[405];
      node522_r = node521_l & pixel[270];
      node522_l = node521_l & ~pixel[270];
      node523_r = node522_l & pixel[189];
      node523_l = node522_l & ~pixel[189];
      node524 = node523_l;
      node525 = node523_r;
      node526_r = node522_r & pixel[595];
      node526_l = node522_r & ~pixel[595];
      node527 = node526_l;
      node528 = node526_r;
      node529_r = node521_r & pixel[232];
      node529_l = node521_r & ~pixel[232];
      node530_r = node529_l & pixel[489];
      node530_l = node529_l & ~pixel[489];
      node531 = node530_l;
      node532 = node530_r;
      node533_r = node529_r & pixel[523];
      node533_l = node529_r & ~pixel[523];
      node534 = node533_l;
      node535 = node533_r;
      node536_r = node520_r & pixel[434];
      node536_l = node520_r & ~pixel[434];
      node537_r = node536_l & pixel[622];
      node537_l = node536_l & ~pixel[622];
      node538_r = node537_l & pixel[493];
      node538_l = node537_l & ~pixel[493];
      node539 = node538_l;
      node540 = node538_r;
      node541 = node537_r;
      node542_r = node536_r & pixel[208];
      node542_l = node536_r & ~pixel[208];
      node543_r = node542_l & pixel[265];
      node543_l = node542_l & ~pixel[265];
      node544 = node543_l;
      node545 = node543_r;
      node546_r = node542_r & pixel[580];
      node546_l = node542_r & ~pixel[580];
      node547 = node546_l;
      node548 = node546_r;
      node549_r = node519_r & pixel[543];
      node549_l = node519_r & ~pixel[543];
      node550_r = node549_l & pixel[346];
      node550_l = node549_l & ~pixel[346];
      node551_r = node550_l & pixel[494];
      node551_l = node550_l & ~pixel[494];
      node552_r = node551_l & pixel[203];
      node552_l = node551_l & ~pixel[203];
      node553 = node552_l;
      node554 = node552_r;
      node555_r = node551_r & pixel[381];
      node555_l = node551_r & ~pixel[381];
      node556 = node555_l;
      node557 = node555_r;
      node558_r = node550_r & pixel[401];
      node558_l = node550_r & ~pixel[401];
      node559_r = node558_l & pixel[269];
      node559_l = node558_l & ~pixel[269];
      node560 = node559_l;
      node561 = node559_r;
      node562_r = node558_r & pixel[596];
      node562_l = node558_r & ~pixel[596];
      node563 = node562_l;
      node564 = node562_r;
      node565_r = node549_r & pixel[293];
      node565_l = node549_r & ~pixel[293];
      node566_r = node565_l & pixel[203];
      node566_l = node565_l & ~pixel[203];
      node567_r = node566_l & pixel[404];
      node567_l = node566_l & ~pixel[404];
      node568 = node567_l;
      node569 = node567_r;
      node570_r = node566_r & pixel[399];
      node570_l = node566_r & ~pixel[399];
      node571 = node570_l;
      node572 = node570_r;
      node573_r = node565_r & pixel[684];
      node573_l = node565_r & ~pixel[684];
      node574_r = node573_l & pixel[639];
      node574_l = node573_l & ~pixel[639];
      node575 = node574_l;
      node576 = node574_r;
      node577_r = node573_r & pixel[380];
      node577_l = node573_r & ~pixel[380];
      node578 = node577_l;
      node579 = node577_r;
      node580_r = node518_r & pixel[469];
      node580_l = node518_r & ~pixel[469];
      node581_r = node580_l & pixel[155];
      node581_l = node580_l & ~pixel[155];
      node582_r = node581_l & pixel[596];
      node582_l = node581_l & ~pixel[596];
      node583_r = node582_l & pixel[211];
      node583_l = node582_l & ~pixel[211];
      node584_r = node583_l & pixel[301];
      node584_l = node583_l & ~pixel[301];
      node585 = node584_l;
      node586 = node584_r;
      node587_r = node583_r & pixel[355];
      node587_l = node583_r & ~pixel[355];
      node588 = node587_l;
      node589 = node587_r;
      node590_r = node582_r & pixel[521];
      node590_l = node582_r & ~pixel[521];
      node591_r = node590_l & pixel[565];
      node591_l = node590_l & ~pixel[565];
      node592 = node591_l;
      node593 = node591_r;
      node594_r = node590_r & pixel[383];
      node594_l = node590_r & ~pixel[383];
      node595 = node594_l;
      node596 = node594_r;
      node597_r = node581_r & pixel[573];
      node597_l = node581_r & ~pixel[573];
      node598_r = node597_l & pixel[685];
      node598_l = node597_l & ~pixel[685];
      node599_r = node598_l & pixel[179];
      node599_l = node598_l & ~pixel[179];
      node600 = node599_l;
      node601 = node599_r;
      node602_r = node598_r & pixel[382];
      node602_l = node598_r & ~pixel[382];
      node603 = node602_l;
      node604 = node602_r;
      node605_r = node597_r & pixel[346];
      node605_l = node597_r & ~pixel[346];
      node606_r = node605_l & pixel[263];
      node606_l = node605_l & ~pixel[263];
      node607 = node606_l;
      node608 = node606_r;
      node609_r = node605_r & pixel[539];
      node609_l = node605_r & ~pixel[539];
      node610 = node609_l;
      node611 = node609_r;
      node612_r = node580_r & pixel[569];
      node612_l = node580_r & ~pixel[569];
      node613_r = node612_l & pixel[719];
      node613_l = node612_l & ~pixel[719];
      node614_r = node613_l & pixel[210];
      node614_l = node613_l & ~pixel[210];
      node615_r = node614_l & pixel[152];
      node615_l = node614_l & ~pixel[152];
      node616 = node615_l;
      node617 = node615_r;
      node618_r = node614_r & pixel[684];
      node618_l = node614_r & ~pixel[684];
      node619 = node618_l;
      node620 = node618_r;
      node621_r = node613_r & pixel[687];
      node621_l = node613_r & ~pixel[687];
      node622_r = node621_l & pixel[472];
      node622_l = node621_l & ~pixel[472];
      node623 = node622_l;
      node624 = node622_r;
      node625_r = node621_r & pixel[631];
      node625_l = node621_r & ~pixel[631];
      node626 = node625_l;
      node627 = node625_r;
      node628_r = node612_r & pixel[347];
      node628_l = node612_r & ~pixel[347];
      node629_r = node628_l & pixel[708];
      node629_l = node628_l & ~pixel[708];
      node630_r = node629_l & pixel[344];
      node630_l = node629_l & ~pixel[344];
      node631 = node630_l;
      node632 = node630_r;
      node633 = node629_r;
      node634_r = node628_r & pixel[244];
      node634_l = node628_r & ~pixel[244];
      node635_r = node634_l & pixel[430];
      node635_l = node634_l & ~pixel[430];
      node636 = node635_l;
      node637 = node635_r;
      node638_r = node634_r & pixel[526];
      node638_l = node634_r & ~pixel[526];
      node639 = node638_l;
      node640 = node638_r;
      node641_r = node397_r & pixel[297];
      node641_l = node397_r & ~pixel[297];
      node642_r = node641_l & pixel[327];
      node642_l = node641_l & ~pixel[327];
      node643_r = node642_l & pixel[487];
      node643_l = node642_l & ~pixel[487];
      node644_r = node643_l & pixel[215];
      node644_l = node643_l & ~pixel[215];
      node645_r = node644_l & pixel[262];
      node645_l = node644_l & ~pixel[262];
      node646_r = node645_l & pixel[206];
      node646_l = node645_l & ~pixel[206];
      node647_r = node646_l & pixel[236];
      node647_l = node646_l & ~pixel[236];
      node648 = node647_l;
      node649 = node647_r;
      node650_r = node646_r & pixel[323];
      node650_l = node646_r & ~pixel[323];
      node651 = node650_l;
      node652 = node650_r;
      node653_r = node645_r & pixel[160];
      node653_l = node645_r & ~pixel[160];
      node654_r = node653_l & pixel[467];
      node654_l = node653_l & ~pixel[467];
      node655 = node654_l;
      node656 = node654_r;
      node657 = node653_r;
      node658_r = node644_r & pixel[356];
      node658_l = node644_r & ~pixel[356];
      node659_r = node658_l & pixel[518];
      node659_l = node658_l & ~pixel[518];
      node660_r = node659_l & pixel[208];
      node660_l = node659_l & ~pixel[208];
      node661 = node660_l;
      node662 = node660_r;
      node663_r = node659_r & pixel[684];
      node663_l = node659_r & ~pixel[684];
      node664 = node663_l;
      node665 = node663_r;
      node666_r = node658_r & pixel[597];
      node666_l = node658_r & ~pixel[597];
      node667_r = node666_l & pixel[539];
      node667_l = node666_l & ~pixel[539];
      node668 = node667_l;
      node669 = node667_r;
      node670_r = node666_r & pixel[124];
      node670_l = node666_r & ~pixel[124];
      node671 = node670_l;
      node672 = node670_r;
      node673_r = node643_r & pixel[655];
      node673_l = node643_r & ~pixel[655];
      node674_r = node673_l & pixel[315];
      node674_l = node673_l & ~pixel[315];
      node675_r = node674_l & pixel[572];
      node675_l = node674_l & ~pixel[572];
      node676_r = node675_l & pixel[215];
      node676_l = node675_l & ~pixel[215];
      node677 = node676_l;
      node678 = node676_r;
      node679_r = node675_r & pixel[656];
      node679_l = node675_r & ~pixel[656];
      node680 = node679_l;
      node681 = node679_r;
      node682_r = node674_r & pixel[211];
      node682_l = node674_r & ~pixel[211];
      node683_r = node682_l & pixel[348];
      node683_l = node682_l & ~pixel[348];
      node684 = node683_l;
      node685 = node683_r;
      node686_r = node682_r & pixel[353];
      node686_l = node682_r & ~pixel[353];
      node687 = node686_l;
      node688 = node686_r;
      node689_r = node673_r & pixel[295];
      node689_l = node673_r & ~pixel[295];
      node690_r = node689_l & pixel[518];
      node690_l = node689_l & ~pixel[518];
      node691_r = node690_l & pixel[298];
      node691_l = node690_l & ~pixel[298];
      node692 = node691_l;
      node693 = node691_r;
      node694_r = node690_r & pixel[493];
      node694_l = node690_r & ~pixel[493];
      node695 = node694_l;
      node696 = node694_r;
      node697_r = node689_r & pixel[323];
      node697_l = node689_r & ~pixel[323];
      node698_r = node697_l & pixel[520];
      node698_l = node697_l & ~pixel[520];
      node699 = node698_l;
      node700 = node698_r;
      node701_r = node697_r & pixel[552];
      node701_l = node697_r & ~pixel[552];
      node702 = node701_l;
      node703 = node701_r;
      node704_r = node642_r & pixel[455];
      node704_l = node642_r & ~pixel[455];
      node705_r = node704_l & pixel[595];
      node705_l = node704_l & ~pixel[595];
      node706_r = node705_l & pixel[658];
      node706_l = node705_l & ~pixel[658];
      node707_r = node706_l & pixel[709];
      node707_l = node706_l & ~pixel[709];
      node708_r = node707_l & pixel[564];
      node708_l = node707_l & ~pixel[564];
      node709 = node708_l;
      node710 = node708_r;
      node711_r = node707_r & pixel[241];
      node711_l = node707_r & ~pixel[241];
      node712 = node711_l;
      node713 = node711_r;
      node714_r = node706_r & pixel[211];
      node714_l = node706_r & ~pixel[211];
      node715_r = node714_l & pixel[516];
      node715_l = node714_l & ~pixel[516];
      node716 = node715_l;
      node717 = node715_r;
      node718_r = node714_r & pixel[402];
      node718_l = node714_r & ~pixel[402];
      node719 = node718_l;
      node720 = node718_r;
      node721_r = node705_r & pixel[379];
      node721_l = node705_r & ~pixel[379];
      node722_r = node721_l & pixel[371];
      node722_l = node721_l & ~pixel[371];
      node723_r = node722_l & pixel[128];
      node723_l = node722_l & ~pixel[128];
      node724 = node723_l;
      node725 = node723_r;
      node726 = node722_r;
      node727_r = node721_r & pixel[320];
      node727_l = node721_r & ~pixel[320];
      node728_r = node727_l & pixel[99];
      node728_l = node727_l & ~pixel[99];
      node729 = node728_l;
      node730 = node728_r;
      node731_r = node727_r & pixel[483];
      node731_l = node727_r & ~pixel[483];
      node732 = node731_l;
      node733 = node731_r;
      node734_r = node704_r & pixel[564];
      node734_l = node704_r & ~pixel[564];
      node735_r = node734_l & pixel[211];
      node735_l = node734_l & ~pixel[211];
      node736_r = node735_l & pixel[213];
      node736_l = node735_l & ~pixel[213];
      node737_r = node736_l & pixel[123];
      node737_l = node736_l & ~pixel[123];
      node738 = node737_l;
      node739 = node737_r;
      node740_r = node736_r & pixel[156];
      node740_l = node736_r & ~pixel[156];
      node741 = node740_l;
      node742 = node740_r;
      node743_r = node735_r & pixel[433];
      node743_l = node735_r & ~pixel[433];
      node744_r = node743_l & pixel[295];
      node744_l = node743_l & ~pixel[295];
      node745 = node744_l;
      node746 = node744_r;
      node747_r = node743_r & pixel[607];
      node747_l = node743_r & ~pixel[607];
      node748 = node747_l;
      node749 = node747_r;
      node750_r = node734_r & pixel[405];
      node750_l = node734_r & ~pixel[405];
      node751 = node750_l;
      node752_r = node750_r & pixel[545];
      node752_l = node750_r & ~pixel[545];
      node753_r = node752_l & pixel[246];
      node753_l = node752_l & ~pixel[246];
      node754 = node753_l;
      node755 = node753_r;
      node756_r = node752_r & pixel[321];
      node756_l = node752_r & ~pixel[321];
      node757 = node756_l;
      node758 = node756_r;
      node759_r = node641_r & pixel[202];
      node759_l = node641_r & ~pixel[202];
      node760_r = node759_l & pixel[157];
      node760_l = node759_l & ~pixel[157];
      node761_r = node760_l & pixel[238];
      node761_l = node760_l & ~pixel[238];
      node762_r = node761_l & pixel[184];
      node762_l = node761_l & ~pixel[184];
      node763_r = node762_l & pixel[403];
      node763_l = node762_l & ~pixel[403];
      node764_r = node763_l & pixel[180];
      node764_l = node763_l & ~pixel[180];
      node765 = node764_l;
      node766 = node764_r;
      node767_r = node763_r & pixel[565];
      node767_l = node763_r & ~pixel[565];
      node768 = node767_l;
      node769 = node767_r;
      node770_r = node762_r & pixel[153];
      node770_l = node762_r & ~pixel[153];
      node771_r = node770_l & pixel[236];
      node771_l = node770_l & ~pixel[236];
      node772 = node771_l;
      node773 = node771_r;
      node774_r = node770_r & pixel[462];
      node774_l = node770_r & ~pixel[462];
      node775 = node774_l;
      node776 = node774_r;
      node777_r = node761_r & pixel[594];
      node777_l = node761_r & ~pixel[594];
      node778_r = node777_l & pixel[149];
      node778_l = node777_l & ~pixel[149];
      node779_r = node778_l & pixel[162];
      node779_l = node778_l & ~pixel[162];
      node780 = node779_l;
      node781 = node779_r;
      node782_r = node778_r & pixel[654];
      node782_l = node778_r & ~pixel[654];
      node783 = node782_l;
      node784 = node782_r;
      node785_r = node777_r & pixel[455];
      node785_l = node777_r & ~pixel[455];
      node786_r = node785_l & pixel[347];
      node786_l = node785_l & ~pixel[347];
      node787 = node786_l;
      node788 = node786_r;
      node789_r = node785_r & pixel[685];
      node789_l = node785_r & ~pixel[685];
      node790 = node789_l;
      node791 = node789_r;
      node792_r = node760_r & pixel[181];
      node792_l = node760_r & ~pixel[181];
      node793_r = node792_l & pixel[519];
      node793_l = node792_l & ~pixel[519];
      node794_r = node793_l & pixel[316];
      node794_l = node793_l & ~pixel[316];
      node795_r = node794_l & pixel[663];
      node795_l = node794_l & ~pixel[663];
      node796 = node795_l;
      node797 = node795_r;
      node798_r = node794_r & pixel[580];
      node798_l = node794_r & ~pixel[580];
      node799 = node798_l;
      node800 = node798_r;
      node801_r = node793_r & pixel[217];
      node801_l = node793_r & ~pixel[217];
      node802_r = node801_l & pixel[598];
      node802_l = node801_l & ~pixel[598];
      node803 = node802_l;
      node804 = node802_r;
      node805_r = node801_r & pixel[513];
      node805_l = node801_r & ~pixel[513];
      node806 = node805_l;
      node807 = node805_r;
      node808_r = node792_r & pixel[622];
      node808_l = node792_r & ~pixel[622];
      node809_r = node808_l & pixel[318];
      node809_l = node808_l & ~pixel[318];
      node810_r = node809_l & pixel[490];
      node810_l = node809_l & ~pixel[490];
      node811 = node810_l;
      node812 = node810_r;
      node813_r = node809_r & pixel[516];
      node813_l = node809_r & ~pixel[516];
      node814 = node813_l;
      node815 = node813_r;
      node816_r = node808_r & pixel[359];
      node816_l = node808_r & ~pixel[359];
      node817_r = node816_l & pixel[316];
      node817_l = node816_l & ~pixel[316];
      node818 = node817_l;
      node819 = node817_r;
      node820_r = node816_r & pixel[649];
      node820_l = node816_r & ~pixel[649];
      node821 = node820_l;
      node822 = node820_r;
      node823_r = node759_r & pixel[368];
      node823_l = node759_r & ~pixel[368];
      node824_r = node823_l & pixel[658];
      node824_l = node823_l & ~pixel[658];
      node825_r = node824_l & pixel[316];
      node825_l = node824_l & ~pixel[316];
      node826_r = node825_l & pixel[177];
      node826_l = node825_l & ~pixel[177];
      node827_r = node826_l & pixel[624];
      node827_l = node826_l & ~pixel[624];
      node828 = node827_l;
      node829 = node827_r;
      node830_r = node826_r & pixel[128];
      node830_l = node826_r & ~pixel[128];
      node831 = node830_l;
      node832 = node830_r;
      node833_r = node825_r & pixel[403];
      node833_l = node825_r & ~pixel[403];
      node834_r = node833_l & pixel[185];
      node834_l = node833_l & ~pixel[185];
      node835 = node834_l;
      node836 = node834_r;
      node837_r = node833_r & pixel[373];
      node837_l = node833_r & ~pixel[373];
      node838 = node837_l;
      node839 = node837_r;
      node840_r = node824_r & pixel[177];
      node840_l = node824_r & ~pixel[177];
      node841_r = node840_l & pixel[355];
      node841_l = node840_l & ~pixel[355];
      node842_r = node841_l & pixel[315];
      node842_l = node841_l & ~pixel[315];
      node843 = node842_l;
      node844 = node842_r;
      node845_r = node841_r & pixel[434];
      node845_l = node841_r & ~pixel[434];
      node846 = node845_l;
      node847 = node845_r;
      node848_r = node840_r & pixel[654];
      node848_l = node840_r & ~pixel[654];
      node849_r = node848_l & pixel[316];
      node849_l = node848_l & ~pixel[316];
      node850 = node849_l;
      node851 = node849_r;
      node852_r = node848_r & pixel[544];
      node852_l = node848_r & ~pixel[544];
      node853 = node852_l;
      node854 = node852_r;
      node855_r = node823_r & pixel[427];
      node855_l = node823_r & ~pixel[427];
      node856_r = node855_l & pixel[689];
      node856_l = node855_l & ~pixel[689];
      node857_r = node856_l & pixel[666];
      node857_l = node856_l & ~pixel[666];
      node858 = node857_l;
      node859 = node857_r;
      node860_r = node856_r & pixel[322];
      node860_l = node856_r & ~pixel[322];
      node861 = node860_l;
      node862 = node860_r;
      node863 = node855_r;
      node864_r = node0_r & pixel[658];
      node864_l = node0_r & ~pixel[658];
      node865_r = node864_l & pixel[319];
      node865_l = node864_l & ~pixel[319];
      node866_r = node865_l & pixel[314];
      node866_l = node865_l & ~pixel[314];
      node867_r = node866_l & pixel[465];
      node867_l = node866_l & ~pixel[465];
      node868_r = node867_l & pixel[155];
      node868_l = node867_l & ~pixel[155];
      node869_r = node868_l & pixel[653];
      node869_l = node868_l & ~pixel[653];
      node870_r = node869_l & pixel[345];
      node870_l = node869_l & ~pixel[345];
      node871_r = node870_l & pixel[208];
      node871_l = node870_l & ~pixel[208];
      node872_r = node871_l & pixel[549];
      node872_l = node871_l & ~pixel[549];
      node873 = node872_l;
      node874 = node872_r;
      node875_r = node871_r & pixel[358];
      node875_l = node871_r & ~pixel[358];
      node876 = node875_l;
      node877 = node875_r;
      node878_r = node870_r & pixel[218];
      node878_l = node870_r & ~pixel[218];
      node879_r = node878_l & pixel[577];
      node879_l = node878_l & ~pixel[577];
      node880 = node879_l;
      node881 = node879_r;
      node882_r = node878_r & pixel[433];
      node882_l = node878_r & ~pixel[433];
      node883 = node882_l;
      node884 = node882_r;
      node885_r = node869_r & pixel[210];
      node885_l = node869_r & ~pixel[210];
      node886_r = node885_l & pixel[438];
      node886_l = node885_l & ~pixel[438];
      node887_r = node886_l & pixel[301];
      node887_l = node886_l & ~pixel[301];
      node888 = node887_l;
      node889 = node887_r;
      node890_r = node886_r & pixel[565];
      node890_l = node886_r & ~pixel[565];
      node891 = node890_l;
      node892 = node890_r;
      node893_r = node885_r & pixel[160];
      node893_l = node885_r & ~pixel[160];
      node894_r = node893_l & pixel[330];
      node894_l = node893_l & ~pixel[330];
      node895 = node894_l;
      node896 = node894_r;
      node897_r = node893_r & pixel[629];
      node897_l = node893_r & ~pixel[629];
      node898 = node897_l;
      node899 = node897_r;
      node900_r = node868_r & pixel[289];
      node900_l = node868_r & ~pixel[289];
      node901_r = node900_l & pixel[207];
      node901_l = node900_l & ~pixel[207];
      node902_r = node901_l & pixel[294];
      node902_l = node901_l & ~pixel[294];
      node903_r = node902_l & pixel[127];
      node903_l = node902_l & ~pixel[127];
      node904 = node903_l;
      node905 = node903_r;
      node906_r = node902_r & pixel[555];
      node906_l = node902_r & ~pixel[555];
      node907 = node906_l;
      node908 = node906_r;
      node909_r = node901_r & pixel[462];
      node909_l = node901_r & ~pixel[462];
      node910_r = node909_l & pixel[485];
      node910_l = node909_l & ~pixel[485];
      node911 = node910_l;
      node912 = node910_r;
      node913_r = node909_r & pixel[320];
      node913_l = node909_r & ~pixel[320];
      node914 = node913_l;
      node915 = node913_r;
      node916_r = node900_r & pixel[441];
      node916_l = node900_r & ~pixel[441];
      node917_r = node916_l & pixel[274];
      node917_l = node916_l & ~pixel[274];
      node918_r = node917_l & pixel[425];
      node918_l = node917_l & ~pixel[425];
      node919 = node918_l;
      node920 = node918_r;
      node921_r = node917_r & pixel[355];
      node921_l = node917_r & ~pixel[355];
      node922 = node921_l;
      node923 = node921_r;
      node924_r = node916_r & pixel[244];
      node924_l = node916_r & ~pixel[244];
      node925_r = node924_l & pixel[427];
      node925_l = node924_l & ~pixel[427];
      node926 = node925_l;
      node927 = node925_r;
      node928_r = node924_r & pixel[491];
      node928_l = node924_r & ~pixel[491];
      node929 = node928_l;
      node930 = node928_r;
      node931_r = node867_r & pixel[316];
      node931_l = node867_r & ~pixel[316];
      node932_r = node931_l & pixel[581];
      node932_l = node931_l & ~pixel[581];
      node933_r = node932_l & pixel[320];
      node933_l = node932_l & ~pixel[320];
      node934_r = node933_l & pixel[709];
      node934_l = node933_l & ~pixel[709];
      node935_r = node934_l & pixel[456];
      node935_l = node934_l & ~pixel[456];
      node936 = node935_l;
      node937 = node935_r;
      node938 = node934_r;
      node939_r = node933_r & pixel[157];
      node939_l = node933_r & ~pixel[157];
      node940_r = node939_l & pixel[330];
      node940_l = node939_l & ~pixel[330];
      node941 = node940_l;
      node942 = node940_r;
      node943_r = node939_r & pixel[154];
      node943_l = node939_r & ~pixel[154];
      node944 = node943_l;
      node945 = node943_r;
      node946_r = node932_r & pixel[258];
      node946_l = node932_r & ~pixel[258];
      node947_r = node946_l & pixel[688];
      node947_l = node946_l & ~pixel[688];
      node948_r = node947_l & pixel[517];
      node948_l = node947_l & ~pixel[517];
      node949 = node948_l;
      node950 = node948_r;
      node951 = node947_r;
      node952_r = node946_r & pixel[353];
      node952_l = node946_r & ~pixel[353];
      node953_r = node952_l & pixel[665];
      node953_l = node952_l & ~pixel[665];
      node954 = node953_l;
      node955 = node953_r;
      node956_r = node952_r & pixel[633];
      node956_l = node952_r & ~pixel[633];
      node957 = node956_l;
      node958 = node956_r;
      node959_r = node931_r & pixel[98];
      node959_l = node931_r & ~pixel[98];
      node960_r = node959_l & pixel[212];
      node960_l = node959_l & ~pixel[212];
      node961_r = node960_l & pixel[400];
      node961_l = node960_l & ~pixel[400];
      node962_r = node961_l & pixel[569];
      node962_l = node961_l & ~pixel[569];
      node963 = node962_l;
      node964 = node962_r;
      node965_r = node961_r & pixel[602];
      node965_l = node961_r & ~pixel[602];
      node966 = node965_l;
      node967 = node965_r;
      node968_r = node960_r & pixel[659];
      node968_l = node960_r & ~pixel[659];
      node969_r = node968_l & pixel[343];
      node969_l = node968_l & ~pixel[343];
      node970 = node969_l;
      node971 = node969_r;
      node972_r = node968_r & pixel[679];
      node972_l = node968_r & ~pixel[679];
      node973 = node972_l;
      node974 = node972_r;
      node975_r = node959_r & pixel[185];
      node975_l = node959_r & ~pixel[185];
      node976 = node975_l;
      node977_r = node975_r & pixel[131];
      node977_l = node975_r & ~pixel[131];
      node978_r = node977_l & pixel[549];
      node978_l = node977_l & ~pixel[549];
      node979 = node978_l;
      node980 = node978_r;
      node981_r = node977_r & pixel[488];
      node981_l = node977_r & ~pixel[488];
      node982 = node981_l;
      node983 = node981_r;
      node984_r = node866_r & pixel[215];
      node984_l = node866_r & ~pixel[215];
      node985_r = node984_l & pixel[270];
      node985_l = node984_l & ~pixel[270];
      node986_r = node985_l & pixel[639];
      node986_l = node985_l & ~pixel[639];
      node987_r = node986_l & pixel[575];
      node987_l = node986_l & ~pixel[575];
      node988_r = node987_l & pixel[328];
      node988_l = node987_l & ~pixel[328];
      node989_r = node988_l & pixel[459];
      node989_l = node988_l & ~pixel[459];
      node990 = node989_l;
      node991 = node989_r;
      node992_r = node988_r & pixel[662];
      node992_l = node988_r & ~pixel[662];
      node993 = node992_l;
      node994 = node992_r;
      node995_r = node987_r & pixel[368];
      node995_l = node987_r & ~pixel[368];
      node996_r = node995_l & pixel[268];
      node996_l = node995_l & ~pixel[268];
      node997 = node996_l;
      node998 = node996_r;
      node999 = node995_r;
      node1000_r = node986_r & pixel[385];
      node1000_l = node986_r & ~pixel[385];
      node1001_r = node1000_l & pixel[230];
      node1001_l = node1000_l & ~pixel[230];
      node1002 = node1001_l;
      node1003 = node1001_r;
      node1004_r = node1000_r & pixel[175];
      node1004_l = node1000_r & ~pixel[175];
      node1005 = node1004_l;
      node1006 = node1004_r;
      node1007_r = node985_r & pixel[406];
      node1007_l = node985_r & ~pixel[406];
      node1008_r = node1007_l & pixel[438];
      node1008_l = node1007_l & ~pixel[438];
      node1009_r = node1008_l & pixel[490];
      node1009_l = node1008_l & ~pixel[490];
      node1010_r = node1009_l & pixel[665];
      node1010_l = node1009_l & ~pixel[665];
      node1011 = node1010_l;
      node1012 = node1010_r;
      node1013_r = node1009_r & pixel[380];
      node1013_l = node1009_r & ~pixel[380];
      node1014 = node1013_l;
      node1015 = node1013_r;
      node1016_r = node1008_r & pixel[630];
      node1016_l = node1008_r & ~pixel[630];
      node1017_r = node1016_l & pixel[370];
      node1017_l = node1016_l & ~pixel[370];
      node1018 = node1017_l;
      node1019 = node1017_r;
      node1020_r = node1016_r & pixel[597];
      node1020_l = node1016_r & ~pixel[597];
      node1021 = node1020_l;
      node1022 = node1020_r;
      node1023_r = node1007_r & pixel[301];
      node1023_l = node1007_r & ~pixel[301];
      node1024_r = node1023_l & pixel[664];
      node1024_l = node1023_l & ~pixel[664];
      node1025_r = node1024_l & pixel[455];
      node1025_l = node1024_l & ~pixel[455];
      node1026 = node1025_l;
      node1027 = node1025_r;
      node1028_r = node1024_r & pixel[375];
      node1028_l = node1024_r & ~pixel[375];
      node1029 = node1028_l;
      node1030 = node1028_r;
      node1031_r = node1023_r & pixel[663];
      node1031_l = node1023_r & ~pixel[663];
      node1032_r = node1031_l & pixel[678];
      node1032_l = node1031_l & ~pixel[678];
      node1033 = node1032_l;
      node1034 = node1032_r;
      node1035_r = node1031_r & pixel[247];
      node1035_l = node1031_r & ~pixel[247];
      node1036 = node1035_l;
      node1037 = node1035_r;
      node1038_r = node984_r & pixel[273];
      node1038_l = node984_r & ~pixel[273];
      node1039_r = node1038_l & pixel[690];
      node1039_l = node1038_l & ~pixel[690];
      node1040_r = node1039_l & pixel[425];
      node1040_l = node1039_l & ~pixel[425];
      node1041_r = node1040_l & pixel[385];
      node1041_l = node1040_l & ~pixel[385];
      node1042_r = node1041_l & pixel[207];
      node1042_l = node1041_l & ~pixel[207];
      node1043 = node1042_l;
      node1044 = node1042_r;
      node1045_r = node1041_r & pixel[519];
      node1045_l = node1041_r & ~pixel[519];
      node1046 = node1045_l;
      node1047 = node1045_r;
      node1048_r = node1040_r & pixel[463];
      node1048_l = node1040_r & ~pixel[463];
      node1049_r = node1048_l & pixel[627];
      node1049_l = node1048_l & ~pixel[627];
      node1050 = node1049_l;
      node1051 = node1049_r;
      node1052_r = node1048_r & pixel[556];
      node1052_l = node1048_r & ~pixel[556];
      node1053 = node1052_l;
      node1054 = node1052_r;
      node1055_r = node1039_r & pixel[202];
      node1055_l = node1039_r & ~pixel[202];
      node1056_r = node1055_l & pixel[522];
      node1056_l = node1055_l & ~pixel[522];
      node1057 = node1056_l;
      node1058 = node1056_r;
      node1059 = node1055_r;
      node1060_r = node1038_r & pixel[184];
      node1060_l = node1038_r & ~pixel[184];
      node1061_r = node1060_l & pixel[470];
      node1061_l = node1060_l & ~pixel[470];
      node1062_r = node1061_l & pixel[486];
      node1062_l = node1061_l & ~pixel[486];
      node1063_r = node1062_l & pixel[663];
      node1063_l = node1062_l & ~pixel[663];
      node1064 = node1063_l;
      node1065 = node1063_r;
      node1066_r = node1062_r & pixel[509];
      node1066_l = node1062_r & ~pixel[509];
      node1067 = node1066_l;
      node1068 = node1066_r;
      node1069_r = node1061_r & pixel[297];
      node1069_l = node1061_r & ~pixel[297];
      node1070_r = node1069_l & pixel[201];
      node1070_l = node1069_l & ~pixel[201];
      node1071 = node1070_l;
      node1072 = node1070_r;
      node1073_r = node1069_r & pixel[452];
      node1073_l = node1069_r & ~pixel[452];
      node1074 = node1073_l;
      node1075 = node1073_r;
      node1076_r = node1060_r & pixel[386];
      node1076_l = node1060_r & ~pixel[386];
      node1077_r = node1076_l & pixel[661];
      node1077_l = node1076_l & ~pixel[661];
      node1078_r = node1077_l & pixel[426];
      node1078_l = node1077_l & ~pixel[426];
      node1079 = node1078_l;
      node1080 = node1078_r;
      node1081_r = node1077_r & pixel[491];
      node1081_l = node1077_r & ~pixel[491];
      node1082 = node1081_l;
      node1083 = node1081_r;
      node1084_r = node1076_r & pixel[599];
      node1084_l = node1076_r & ~pixel[599];
      node1085_r = node1084_l & pixel[496];
      node1085_l = node1084_l & ~pixel[496];
      node1086 = node1085_l;
      node1087 = node1085_r;
      node1088_r = node1084_r & pixel[343];
      node1088_l = node1084_r & ~pixel[343];
      node1089 = node1088_l;
      node1090 = node1088_r;
      node1091_r = node865_r & pixel[101];
      node1091_l = node865_r & ~pixel[101];
      node1092_r = node1091_l & pixel[216];
      node1092_l = node1091_l & ~pixel[216];
      node1093_r = node1092_l & pixel[246];
      node1093_l = node1092_l & ~pixel[246];
      node1094_r = node1093_l & pixel[300];
      node1094_l = node1093_l & ~pixel[300];
      node1095_r = node1094_l & pixel[325];
      node1095_l = node1094_l & ~pixel[325];
      node1096_r = node1095_l & pixel[429];
      node1096_l = node1095_l & ~pixel[429];
      node1097_r = node1096_l & pixel[461];
      node1097_l = node1096_l & ~pixel[461];
      node1098 = node1097_l;
      node1099 = node1097_r;
      node1100_r = node1096_r & pixel[92];
      node1100_l = node1096_r & ~pixel[92];
      node1101 = node1100_l;
      node1102 = node1100_r;
      node1103_r = node1095_r & pixel[69];
      node1103_l = node1095_r & ~pixel[69];
      node1104_r = node1103_l & pixel[296];
      node1104_l = node1103_l & ~pixel[296];
      node1105 = node1104_l;
      node1106 = node1104_r;
      node1107 = node1103_r;
      node1108_r = node1094_r & pixel[380];
      node1108_l = node1094_r & ~pixel[380];
      node1109_r = node1108_l & pixel[404];
      node1109_l = node1108_l & ~pixel[404];
      node1110_r = node1109_l & pixel[241];
      node1110_l = node1109_l & ~pixel[241];
      node1111 = node1110_l;
      node1112 = node1110_r;
      node1113_r = node1109_r & pixel[157];
      node1113_l = node1109_r & ~pixel[157];
      node1114 = node1113_l;
      node1115 = node1113_r;
      node1116_r = node1108_r & pixel[243];
      node1116_l = node1108_r & ~pixel[243];
      node1117_r = node1116_l & pixel[124];
      node1117_l = node1116_l & ~pixel[124];
      node1118 = node1117_l;
      node1119 = node1117_r;
      node1120_r = node1116_r & pixel[601];
      node1120_l = node1116_r & ~pixel[601];
      node1121 = node1120_l;
      node1122 = node1120_r;
      node1123_r = node1093_r & pixel[294];
      node1123_l = node1093_r & ~pixel[294];
      node1124_r = node1123_l & pixel[371];
      node1124_l = node1123_l & ~pixel[371];
      node1125_r = node1124_l & pixel[401];
      node1125_l = node1124_l & ~pixel[401];
      node1126_r = node1125_l & pixel[509];
      node1126_l = node1125_l & ~pixel[509];
      node1127 = node1126_l;
      node1128 = node1126_r;
      node1129_r = node1125_r & pixel[184];
      node1129_l = node1125_r & ~pixel[184];
      node1130 = node1129_l;
      node1131 = node1129_r;
      node1132_r = node1124_r & pixel[160];
      node1132_l = node1124_r & ~pixel[160];
      node1133_r = node1132_l & pixel[210];
      node1133_l = node1132_l & ~pixel[210];
      node1134 = node1133_l;
      node1135 = node1133_r;
      node1136 = node1132_r;
      node1137_r = node1123_r & pixel[383];
      node1137_l = node1123_r & ~pixel[383];
      node1138_r = node1137_l & pixel[654];
      node1138_l = node1137_l & ~pixel[654];
      node1139_r = node1138_l & pixel[499];
      node1139_l = node1138_l & ~pixel[499];
      node1140 = node1139_l;
      node1141 = node1139_r;
      node1142_r = node1138_r & pixel[488];
      node1142_l = node1138_r & ~pixel[488];
      node1143 = node1142_l;
      node1144 = node1142_r;
      node1145_r = node1137_r & pixel[242];
      node1145_l = node1137_r & ~pixel[242];
      node1146_r = node1145_l & pixel[300];
      node1146_l = node1145_l & ~pixel[300];
      node1147 = node1146_l;
      node1148 = node1146_r;
      node1149_r = node1145_r & pixel[511];
      node1149_l = node1145_r & ~pixel[511];
      node1150 = node1149_l;
      node1151 = node1149_r;
      node1152_r = node1092_r & pixel[487];
      node1152_l = node1092_r & ~pixel[487];
      node1153_r = node1152_l & pixel[386];
      node1153_l = node1152_l & ~pixel[386];
      node1154_r = node1153_l & pixel[326];
      node1154_l = node1153_l & ~pixel[326];
      node1155_r = node1154_l & pixel[413];
      node1155_l = node1154_l & ~pixel[413];
      node1156_r = node1155_l & pixel[412];
      node1156_l = node1155_l & ~pixel[412];
      node1157 = node1156_l;
      node1158 = node1156_r;
      node1159_r = node1155_r & pixel[160];
      node1159_l = node1155_r & ~pixel[160];
      node1160 = node1159_l;
      node1161 = node1159_r;
      node1162_r = node1154_r & pixel[536];
      node1162_l = node1154_r & ~pixel[536];
      node1163_r = node1162_l & pixel[485];
      node1163_l = node1162_l & ~pixel[485];
      node1164 = node1163_l;
      node1165 = node1163_r;
      node1166_r = node1162_r & pixel[299];
      node1166_l = node1162_r & ~pixel[299];
      node1167 = node1166_l;
      node1168 = node1166_r;
      node1169_r = node1153_r & pixel[407];
      node1169_l = node1153_r & ~pixel[407];
      node1170_r = node1169_l & pixel[203];
      node1170_l = node1169_l & ~pixel[203];
      node1171_r = node1170_l & pixel[573];
      node1171_l = node1170_l & ~pixel[573];
      node1172 = node1171_l;
      node1173 = node1171_r;
      node1174_r = node1170_r & pixel[554];
      node1174_l = node1170_r & ~pixel[554];
      node1175 = node1174_l;
      node1176 = node1174_r;
      node1177_r = node1169_r & pixel[292];
      node1177_l = node1169_r & ~pixel[292];
      node1178 = node1177_l;
      node1179_r = node1177_r & pixel[213];
      node1179_l = node1177_r & ~pixel[213];
      node1180 = node1179_l;
      node1181 = node1179_r;
      node1182_r = node1152_r & pixel[456];
      node1182_l = node1152_r & ~pixel[456];
      node1183_r = node1182_l & pixel[656];
      node1183_l = node1182_l & ~pixel[656];
      node1184_r = node1183_l & pixel[299];
      node1184_l = node1183_l & ~pixel[299];
      node1185_r = node1184_l & pixel[455];
      node1185_l = node1184_l & ~pixel[455];
      node1186 = node1185_l;
      node1187 = node1185_r;
      node1188_r = node1184_r & pixel[707];
      node1188_l = node1184_r & ~pixel[707];
      node1189 = node1188_l;
      node1190 = node1188_r;
      node1191_r = node1183_r & pixel[316];
      node1191_l = node1183_r & ~pixel[316];
      node1192_r = node1191_l & pixel[715];
      node1192_l = node1191_l & ~pixel[715];
      node1193 = node1192_l;
      node1194 = node1192_r;
      node1195_r = node1191_r & pixel[184];
      node1195_l = node1191_r & ~pixel[184];
      node1196 = node1195_l;
      node1197 = node1195_r;
      node1198_r = node1182_r & pixel[374];
      node1198_l = node1182_r & ~pixel[374];
      node1199_r = node1198_l & pixel[212];
      node1199_l = node1198_l & ~pixel[212];
      node1200_r = node1199_l & pixel[129];
      node1200_l = node1199_l & ~pixel[129];
      node1201 = node1200_l;
      node1202 = node1200_r;
      node1203_r = node1199_r & pixel[657];
      node1203_l = node1199_r & ~pixel[657];
      node1204 = node1203_l;
      node1205 = node1203_r;
      node1206_r = node1198_r & pixel[183];
      node1206_l = node1198_r & ~pixel[183];
      node1207_r = node1206_l & pixel[318];
      node1207_l = node1206_l & ~pixel[318];
      node1208 = node1207_l;
      node1209 = node1207_r;
      node1210_r = node1206_r & pixel[105];
      node1210_l = node1206_r & ~pixel[105];
      node1211 = node1210_l;
      node1212 = node1210_r;
      node1213_r = node1091_r & pixel[623];
      node1213_l = node1091_r & ~pixel[623];
      node1214_r = node1213_l & pixel[124];
      node1214_l = node1213_l & ~pixel[124];
      node1215_r = node1214_l & pixel[537];
      node1215_l = node1214_l & ~pixel[537];
      node1216_r = node1215_l & pixel[245];
      node1216_l = node1215_l & ~pixel[245];
      node1217_r = node1216_l & pixel[244];
      node1217_l = node1216_l & ~pixel[244];
      node1218_r = node1217_l & pixel[150];
      node1218_l = node1217_l & ~pixel[150];
      node1219 = node1218_l;
      node1220 = node1218_r;
      node1221_r = node1217_r & pixel[435];
      node1221_l = node1217_r & ~pixel[435];
      node1222 = node1221_l;
      node1223 = node1221_r;
      node1224_r = node1216_r & pixel[463];
      node1224_l = node1216_r & ~pixel[463];
      node1225_r = node1224_l & pixel[290];
      node1225_l = node1224_l & ~pixel[290];
      node1226 = node1225_l;
      node1227 = node1225_r;
      node1228 = node1224_r;
      node1229_r = node1215_r & pixel[442];
      node1229_l = node1215_r & ~pixel[442];
      node1230_r = node1229_l & pixel[271];
      node1230_l = node1229_l & ~pixel[271];
      node1231_r = node1230_l & pixel[102];
      node1231_l = node1230_l & ~pixel[102];
      node1232 = node1231_l;
      node1233 = node1231_r;
      node1234_r = node1230_r & pixel[622];
      node1234_l = node1230_r & ~pixel[622];
      node1235 = node1234_l;
      node1236 = node1234_r;
      node1237_r = node1229_r & pixel[368];
      node1237_l = node1229_r & ~pixel[368];
      node1238_r = node1237_l & pixel[413];
      node1238_l = node1237_l & ~pixel[413];
      node1239 = node1238_l;
      node1240 = node1238_r;
      node1241 = node1237_r;
      node1242_r = node1214_r & pixel[400];
      node1242_l = node1214_r & ~pixel[400];
      node1243_r = node1242_l & pixel[235];
      node1243_l = node1242_l & ~pixel[235];
      node1244_r = node1243_l & pixel[238];
      node1244_l = node1243_l & ~pixel[238];
      node1245_r = node1244_l & pixel[522];
      node1245_l = node1244_l & ~pixel[522];
      node1246 = node1245_l;
      node1247 = node1245_r;
      node1248_r = node1244_r & pixel[158];
      node1248_l = node1244_r & ~pixel[158];
      node1249 = node1248_l;
      node1250 = node1248_r;
      node1251_r = node1243_r & pixel[467];
      node1251_l = node1243_r & ~pixel[467];
      node1252_r = node1251_l & pixel[470];
      node1252_l = node1251_l & ~pixel[470];
      node1253 = node1252_l;
      node1254 = node1252_r;
      node1255_r = node1251_r & pixel[492];
      node1255_l = node1251_r & ~pixel[492];
      node1256 = node1255_l;
      node1257 = node1255_r;
      node1258_r = node1242_r & pixel[290];
      node1258_l = node1242_r & ~pixel[290];
      node1259_r = node1258_l & pixel[370];
      node1259_l = node1258_l & ~pixel[370];
      node1260_r = node1259_l & pixel[517];
      node1260_l = node1259_l & ~pixel[517];
      node1261 = node1260_l;
      node1262 = node1260_r;
      node1263 = node1259_r;
      node1264_r = node1258_r & pixel[434];
      node1264_l = node1258_r & ~pixel[434];
      node1265_r = node1264_l & pixel[410];
      node1265_l = node1264_l & ~pixel[410];
      node1266 = node1265_l;
      node1267 = node1265_r;
      node1268 = node1264_r;
      node1269_r = node1213_r & pixel[593];
      node1269_l = node1213_r & ~pixel[593];
      node1270_r = node1269_l & pixel[429];
      node1270_l = node1269_l & ~pixel[429];
      node1271_r = node1270_l & pixel[628];
      node1271_l = node1270_l & ~pixel[628];
      node1272_r = node1271_l & pixel[550];
      node1272_l = node1271_l & ~pixel[550];
      node1273 = node1272_l;
      node1274_r = node1272_r & pixel[411];
      node1274_l = node1272_r & ~pixel[411];
      node1275 = node1274_l;
      node1276 = node1274_r;
      node1277_r = node1271_r & pixel[261];
      node1277_l = node1271_r & ~pixel[261];
      node1278 = node1277_l;
      node1279_r = node1277_r & pixel[455];
      node1279_l = node1277_r & ~pixel[455];
      node1280 = node1279_l;
      node1281 = node1279_r;
      node1282_r = node1270_r & pixel[437];
      node1282_l = node1270_r & ~pixel[437];
      node1283_r = node1282_l & pixel[244];
      node1283_l = node1282_l & ~pixel[244];
      node1284 = node1283_l;
      node1285 = node1283_r;
      node1286_r = node1282_r & pixel[298];
      node1286_l = node1282_r & ~pixel[298];
      node1287 = node1286_l;
      node1288_r = node1286_r & pixel[331];
      node1288_l = node1286_r & ~pixel[331];
      node1289 = node1288_l;
      node1290 = node1288_r;
      node1291_r = node1269_r & pixel[324];
      node1291_l = node1269_r & ~pixel[324];
      node1292_r = node1291_l & pixel[326];
      node1292_l = node1291_l & ~pixel[326];
      node1293_r = node1292_l & pixel[428];
      node1293_l = node1292_l & ~pixel[428];
      node1294_r = node1293_l & pixel[262];
      node1294_l = node1293_l & ~pixel[262];
      node1295 = node1294_l;
      node1296 = node1294_r;
      node1297_r = node1293_r & pixel[213];
      node1297_l = node1293_r & ~pixel[213];
      node1298 = node1297_l;
      node1299 = node1297_r;
      node1300_r = node1292_r & pixel[408];
      node1300_l = node1292_r & ~pixel[408];
      node1301 = node1300_l;
      node1302 = node1300_r;
      node1303_r = node1291_r & pixel[497];
      node1303_l = node1291_r & ~pixel[497];
      node1304_r = node1303_l & pixel[540];
      node1304_l = node1303_l & ~pixel[540];
      node1305 = node1304_l;
      node1306 = node1304_r;
      node1307_r = node1303_r & pixel[507];
      node1307_l = node1303_r & ~pixel[507];
      node1308_r = node1307_l & pixel[104];
      node1308_l = node1307_l & ~pixel[104];
      node1309 = node1308_l;
      node1310 = node1308_r;
      node1311 = node1307_r;
      node1312_r = node864_r & pixel[377];
      node1312_l = node864_r & ~pixel[377];
      node1313_r = node1312_l & pixel[463];
      node1313_l = node1312_l & ~pixel[463];
      node1314_r = node1313_l & pixel[214];
      node1314_l = node1313_l & ~pixel[214];
      node1315_r = node1314_l & pixel[484];
      node1315_l = node1314_l & ~pixel[484];
      node1316_r = node1315_l & pixel[350];
      node1316_l = node1315_l & ~pixel[350];
      node1317_r = node1316_l & pixel[407];
      node1317_l = node1316_l & ~pixel[407];
      node1318_r = node1317_l & pixel[433];
      node1318_l = node1317_l & ~pixel[433];
      node1319_r = node1318_l & pixel[149];
      node1319_l = node1318_l & ~pixel[149];
      node1320 = node1319_l;
      node1321 = node1319_r;
      node1322 = node1318_r;
      node1323_r = node1317_r & pixel[663];
      node1323_l = node1317_r & ~pixel[663];
      node1324_r = node1323_l & pixel[500];
      node1324_l = node1323_l & ~pixel[500];
      node1325 = node1324_l;
      node1326 = node1324_r;
      node1327 = node1323_r;
      node1328_r = node1316_r & pixel[440];
      node1328_l = node1316_r & ~pixel[440];
      node1329_r = node1328_l & pixel[432];
      node1329_l = node1328_l & ~pixel[432];
      node1330_r = node1329_l & pixel[185];
      node1330_l = node1329_l & ~pixel[185];
      node1331 = node1330_l;
      node1332 = node1330_r;
      node1333 = node1329_r;
      node1334_r = node1328_r & pixel[331];
      node1334_l = node1328_r & ~pixel[331];
      node1335_r = node1334_l & pixel[128];
      node1335_l = node1334_l & ~pixel[128];
      node1336 = node1335_l;
      node1337 = node1335_r;
      node1338 = node1334_r;
      node1339_r = node1315_r & pixel[147];
      node1339_l = node1315_r & ~pixel[147];
      node1340_r = node1339_l & pixel[378];
      node1340_l = node1339_l & ~pixel[378];
      node1341_r = node1340_l & pixel[372];
      node1341_l = node1340_l & ~pixel[372];
      node1342_r = node1341_l & pixel[295];
      node1342_l = node1341_l & ~pixel[295];
      node1343 = node1342_l;
      node1344 = node1342_r;
      node1345_r = node1341_r & pixel[657];
      node1345_l = node1341_r & ~pixel[657];
      node1346 = node1345_l;
      node1347 = node1345_r;
      node1348_r = node1340_r & pixel[263];
      node1348_l = node1340_r & ~pixel[263];
      node1349_r = node1348_l & pixel[429];
      node1349_l = node1348_l & ~pixel[429];
      node1350 = node1349_l;
      node1351 = node1349_r;
      node1352_r = node1348_r & pixel[486];
      node1352_l = node1348_r & ~pixel[486];
      node1353 = node1352_l;
      node1354 = node1352_r;
      node1355_r = node1339_r & pixel[483];
      node1355_l = node1339_r & ~pixel[483];
      node1356_r = node1355_l & pixel[288];
      node1356_l = node1355_l & ~pixel[288];
      node1357_r = node1356_l & pixel[465];
      node1357_l = node1356_l & ~pixel[465];
      node1358 = node1357_l;
      node1359 = node1357_r;
      node1360 = node1356_r;
      node1361_r = node1355_r & pixel[293];
      node1361_l = node1355_r & ~pixel[293];
      node1362 = node1361_l;
      node1363_r = node1361_r & pixel[472];
      node1363_l = node1361_r & ~pixel[472];
      node1364 = node1363_l;
      node1365 = node1363_r;
      node1366_r = node1314_r & pixel[433];
      node1366_l = node1314_r & ~pixel[433];
      node1367_r = node1366_l & pixel[349];
      node1367_l = node1366_l & ~pixel[349];
      node1368_r = node1367_l & pixel[382];
      node1368_l = node1367_l & ~pixel[382];
      node1369_r = node1368_l & pixel[434];
      node1369_l = node1368_l & ~pixel[434];
      node1370_r = node1369_l & pixel[488];
      node1370_l = node1369_l & ~pixel[488];
      node1371 = node1370_l;
      node1372 = node1370_r;
      node1373 = node1369_r;
      node1374_r = node1368_r & pixel[351];
      node1374_l = node1368_r & ~pixel[351];
      node1375_r = node1374_l & pixel[154];
      node1375_l = node1374_l & ~pixel[154];
      node1376 = node1375_l;
      node1377 = node1375_r;
      node1378_r = node1374_r & pixel[384];
      node1378_l = node1374_r & ~pixel[384];
      node1379 = node1378_l;
      node1380 = node1378_r;
      node1381_r = node1367_r & pixel[151];
      node1381_l = node1367_r & ~pixel[151];
      node1382_r = node1381_l & pixel[242];
      node1382_l = node1381_l & ~pixel[242];
      node1383_r = node1382_l & pixel[574];
      node1383_l = node1382_l & ~pixel[574];
      node1384 = node1383_l;
      node1385 = node1383_r;
      node1386_r = node1382_r & pixel[328];
      node1386_l = node1382_r & ~pixel[328];
      node1387 = node1386_l;
      node1388 = node1386_r;
      node1389_r = node1381_r & pixel[216];
      node1389_l = node1381_r & ~pixel[216];
      node1390_r = node1389_l & pixel[268];
      node1390_l = node1389_l & ~pixel[268];
      node1391 = node1390_l;
      node1392 = node1390_r;
      node1393_r = node1389_r & pixel[330];
      node1393_l = node1389_r & ~pixel[330];
      node1394 = node1393_l;
      node1395 = node1393_r;
      node1396_r = node1366_r & pixel[633];
      node1396_l = node1366_r & ~pixel[633];
      node1397_r = node1396_l & pixel[221];
      node1397_l = node1396_l & ~pixel[221];
      node1398_r = node1397_l & pixel[453];
      node1398_l = node1397_l & ~pixel[453];
      node1399_r = node1398_l & pixel[689];
      node1399_l = node1398_l & ~pixel[689];
      node1400 = node1399_l;
      node1401 = node1399_r;
      node1402 = node1398_r;
      node1403_r = node1397_r & pixel[660];
      node1403_l = node1397_r & ~pixel[660];
      node1404 = node1403_l;
      node1405 = node1403_r;
      node1406_r = node1396_r & pixel[401];
      node1406_l = node1396_r & ~pixel[401];
      node1407_r = node1406_l & pixel[289];
      node1407_l = node1406_l & ~pixel[289];
      node1408_r = node1407_l & pixel[376];
      node1408_l = node1407_l & ~pixel[376];
      node1409 = node1408_l;
      node1410 = node1408_r;
      node1411_r = node1407_r & pixel[330];
      node1411_l = node1407_r & ~pixel[330];
      node1412 = node1411_l;
      node1413 = node1411_r;
      node1414_r = node1406_r & pixel[356];
      node1414_l = node1406_r & ~pixel[356];
      node1415 = node1414_l;
      node1416 = node1414_r;
      node1417_r = node1313_r & pixel[402];
      node1417_l = node1313_r & ~pixel[402];
      node1418_r = node1417_l & pixel[634];
      node1418_l = node1417_l & ~pixel[634];
      node1419_r = node1418_l & pixel[427];
      node1419_l = node1418_l & ~pixel[427];
      node1420_r = node1419_l & pixel[352];
      node1420_l = node1419_l & ~pixel[352];
      node1421_r = node1420_l & pixel[714];
      node1421_l = node1420_l & ~pixel[714];
      node1422_r = node1421_l & pixel[466];
      node1422_l = node1421_l & ~pixel[466];
      node1423 = node1422_l;
      node1424 = node1422_r;
      node1425_r = node1421_r & pixel[712];
      node1425_l = node1421_r & ~pixel[712];
      node1426 = node1425_l;
      node1427 = node1425_r;
      node1428_r = node1420_r & pixel[682];
      node1428_l = node1420_r & ~pixel[682];
      node1429_r = node1428_l & pixel[713];
      node1429_l = node1428_l & ~pixel[713];
      node1430 = node1429_l;
      node1431 = node1429_r;
      node1432_r = node1428_r & pixel[606];
      node1432_l = node1428_r & ~pixel[606];
      node1433 = node1432_l;
      node1434 = node1432_r;
      node1435_r = node1419_r & pixel[713];
      node1435_l = node1419_r & ~pixel[713];
      node1436_r = node1435_l & pixel[211];
      node1436_l = node1435_l & ~pixel[211];
      node1437_r = node1436_l & pixel[428];
      node1437_l = node1436_l & ~pixel[428];
      node1438 = node1437_l;
      node1439 = node1437_r;
      node1440_r = node1436_r & pixel[384];
      node1440_l = node1436_r & ~pixel[384];
      node1441 = node1440_l;
      node1442 = node1440_r;
      node1443_r = node1435_r & pixel[625];
      node1443_l = node1435_r & ~pixel[625];
      node1444_r = node1443_l & pixel[204];
      node1444_l = node1443_l & ~pixel[204];
      node1445 = node1444_l;
      node1446 = node1444_r;
      node1447 = node1443_r;
      node1448_r = node1418_r & pixel[330];
      node1448_l = node1418_r & ~pixel[330];
      node1449_r = node1448_l & pixel[345];
      node1449_l = node1448_l & ~pixel[345];
      node1450_r = node1449_l & pixel[497];
      node1450_l = node1449_l & ~pixel[497];
      node1451_r = node1450_l & pixel[152];
      node1451_l = node1450_l & ~pixel[152];
      node1452 = node1451_l;
      node1453 = node1451_r;
      node1454_r = node1450_r & pixel[427];
      node1454_l = node1450_r & ~pixel[427];
      node1455 = node1454_l;
      node1456 = node1454_r;
      node1457_r = node1449_r & pixel[485];
      node1457_l = node1449_r & ~pixel[485];
      node1458 = node1457_l;
      node1459_r = node1457_r & pixel[511];
      node1459_l = node1457_r & ~pixel[511];
      node1460 = node1459_l;
      node1461 = node1459_r;
      node1462_r = node1448_r & pixel[655];
      node1462_l = node1448_r & ~pixel[655];
      node1463_r = node1462_l & pixel[325];
      node1463_l = node1462_l & ~pixel[325];
      node1464_r = node1463_l & pixel[236];
      node1464_l = node1463_l & ~pixel[236];
      node1465 = node1464_l;
      node1466 = node1464_r;
      node1467 = node1463_r;
      node1468_r = node1462_r & pixel[371];
      node1468_l = node1462_r & ~pixel[371];
      node1469 = node1468_l;
      node1470_r = node1468_r & pixel[604];
      node1470_l = node1468_r & ~pixel[604];
      node1471 = node1470_l;
      node1472 = node1470_r;
      node1473_r = node1417_r & pixel[403];
      node1473_l = node1417_r & ~pixel[403];
      node1474_r = node1473_l & pixel[547];
      node1474_l = node1473_l & ~pixel[547];
      node1475_r = node1474_l & pixel[683];
      node1475_l = node1474_l & ~pixel[683];
      node1476_r = node1475_l & pixel[357];
      node1476_l = node1475_l & ~pixel[357];
      node1477_r = node1476_l & pixel[204];
      node1477_l = node1476_l & ~pixel[204];
      node1478 = node1477_l;
      node1479 = node1477_r;
      node1480 = node1476_r;
      node1481_r = node1475_r & pixel[545];
      node1481_l = node1475_r & ~pixel[545];
      node1482 = node1481_l;
      node1483 = node1481_r;
      node1484_r = node1474_r & pixel[185];
      node1484_l = node1474_r & ~pixel[185];
      node1485_r = node1484_l & pixel[680];
      node1485_l = node1484_l & ~pixel[680];
      node1486 = node1485_l;
      node1487 = node1485_r;
      node1488_r = node1484_r & pixel[653];
      node1488_l = node1484_r & ~pixel[653];
      node1489_r = node1488_l & pixel[442];
      node1489_l = node1488_l & ~pixel[442];
      node1490 = node1489_l;
      node1491 = node1489_r;
      node1492_r = node1488_r & pixel[347];
      node1492_l = node1488_r & ~pixel[347];
      node1493 = node1492_l;
      node1494 = node1492_r;
      node1495_r = node1473_r & pixel[348];
      node1495_l = node1473_r & ~pixel[348];
      node1496_r = node1495_l & pixel[514];
      node1496_l = node1495_l & ~pixel[514];
      node1497_r = node1496_l & pixel[412];
      node1497_l = node1496_l & ~pixel[412];
      node1498_r = node1497_l & pixel[344];
      node1498_l = node1497_l & ~pixel[344];
      node1499 = node1498_l;
      node1500 = node1498_r;
      node1501_r = node1497_r & pixel[173];
      node1501_l = node1497_r & ~pixel[173];
      node1502 = node1501_l;
      node1503 = node1501_r;
      node1504_r = node1496_r & pixel[654];
      node1504_l = node1496_r & ~pixel[654];
      node1505_r = node1504_l & pixel[318];
      node1505_l = node1504_l & ~pixel[318];
      node1506 = node1505_l;
      node1507 = node1505_r;
      node1508_r = node1504_r & pixel[556];
      node1508_l = node1504_r & ~pixel[556];
      node1509 = node1508_l;
      node1510 = node1508_r;
      node1511_r = node1495_r & pixel[465];
      node1511_l = node1495_r & ~pixel[465];
      node1512_r = node1511_l & pixel[680];
      node1512_l = node1511_l & ~pixel[680];
      node1513_r = node1512_l & pixel[483];
      node1513_l = node1512_l & ~pixel[483];
      node1514 = node1513_l;
      node1515 = node1513_r;
      node1516_r = node1512_r & pixel[457];
      node1516_l = node1512_r & ~pixel[457];
      node1517 = node1516_l;
      node1518 = node1516_r;
      node1519_r = node1511_r & pixel[713];
      node1519_l = node1511_r & ~pixel[713];
      node1520_r = node1519_l & pixel[352];
      node1520_l = node1519_l & ~pixel[352];
      node1521 = node1520_l;
      node1522 = node1520_r;
      node1523 = node1519_r;
      node1524_r = node1312_r & pixel[272];
      node1524_l = node1312_r & ~pixel[272];
      node1525_r = node1524_l & pixel[290];
      node1525_l = node1524_l & ~pixel[290];
      node1526_r = node1525_l & pixel[515];
      node1526_l = node1525_l & ~pixel[515];
      node1527_r = node1526_l & pixel[292];
      node1527_l = node1526_l & ~pixel[292];
      node1528_r = node1527_l & pixel[296];
      node1528_l = node1527_l & ~pixel[296];
      node1529_r = node1528_l & pixel[373];
      node1529_l = node1528_l & ~pixel[373];
      node1530_r = node1529_l & pixel[245];
      node1530_l = node1529_l & ~pixel[245];
      node1531 = node1530_l;
      node1532 = node1530_r;
      node1533_r = node1529_r & pixel[204];
      node1533_l = node1529_r & ~pixel[204];
      node1534 = node1533_l;
      node1535 = node1533_r;
      node1536_r = node1528_r & pixel[611];
      node1536_l = node1528_r & ~pixel[611];
      node1537_r = node1536_l & pixel[350];
      node1537_l = node1536_l & ~pixel[350];
      node1538 = node1537_l;
      node1539 = node1537_r;
      node1540_r = node1536_r & pixel[571];
      node1540_l = node1536_r & ~pixel[571];
      node1541 = node1540_l;
      node1542 = node1540_r;
      node1543_r = node1527_r & pixel[148];
      node1543_l = node1527_r & ~pixel[148];
      node1544_r = node1543_l & pixel[164];
      node1544_l = node1543_l & ~pixel[164];
      node1545_r = node1544_l & pixel[177];
      node1545_l = node1544_l & ~pixel[177];
      node1546 = node1545_l;
      node1547 = node1545_r;
      node1548_r = node1544_r & pixel[519];
      node1548_l = node1544_r & ~pixel[519];
      node1549 = node1548_l;
      node1550 = node1548_r;
      node1551_r = node1543_r & pixel[427];
      node1551_l = node1543_r & ~pixel[427];
      node1552_r = node1551_l & pixel[689];
      node1552_l = node1551_l & ~pixel[689];
      node1553 = node1552_l;
      node1554 = node1552_r;
      node1555_r = node1551_r & pixel[295];
      node1555_l = node1551_r & ~pixel[295];
      node1556 = node1555_l;
      node1557 = node1555_r;
      node1558_r = node1526_r & pixel[438];
      node1558_l = node1526_r & ~pixel[438];
      node1559_r = node1558_l & pixel[636];
      node1559_l = node1558_l & ~pixel[636];
      node1560_r = node1559_l & pixel[150];
      node1560_l = node1559_l & ~pixel[150];
      node1561_r = node1560_l & pixel[401];
      node1561_l = node1560_l & ~pixel[401];
      node1562 = node1561_l;
      node1563 = node1561_r;
      node1564_r = node1560_r & pixel[258];
      node1564_l = node1560_r & ~pixel[258];
      node1565 = node1564_l;
      node1566 = node1564_r;
      node1567_r = node1559_r & pixel[400];
      node1567_l = node1559_r & ~pixel[400];
      node1568_r = node1567_l & pixel[289];
      node1568_l = node1567_l & ~pixel[289];
      node1569 = node1568_l;
      node1570 = node1568_r;
      node1571_r = node1567_r & pixel[230];
      node1571_l = node1567_r & ~pixel[230];
      node1572 = node1571_l;
      node1573 = node1571_r;
      node1574_r = node1558_r & pixel[122];
      node1574_l = node1558_r & ~pixel[122];
      node1575_r = node1574_l & pixel[180];
      node1575_l = node1574_l & ~pixel[180];
      node1576_r = node1575_l & pixel[349];
      node1576_l = node1575_l & ~pixel[349];
      node1577 = node1576_l;
      node1578 = node1576_r;
      node1579_r = node1575_r & pixel[459];
      node1579_l = node1575_r & ~pixel[459];
      node1580 = node1579_l;
      node1581 = node1579_r;
      node1582_r = node1574_r & pixel[555];
      node1582_l = node1574_r & ~pixel[555];
      node1583_r = node1582_l & pixel[120];
      node1583_l = node1582_l & ~pixel[120];
      node1584 = node1583_l;
      node1585 = node1583_r;
      node1586_r = node1582_r & pixel[519];
      node1586_l = node1582_r & ~pixel[519];
      node1587 = node1586_l;
      node1588 = node1586_r;
      node1589_r = node1525_r & pixel[298];
      node1589_l = node1525_r & ~pixel[298];
      node1590_r = node1589_l & pixel[328];
      node1590_l = node1589_l & ~pixel[328];
      node1591_r = node1590_l & pixel[158];
      node1591_l = node1590_l & ~pixel[158];
      node1592_r = node1591_l & pixel[322];
      node1592_l = node1591_l & ~pixel[322];
      node1593_r = node1592_l & pixel[551];
      node1593_l = node1592_l & ~pixel[551];
      node1594 = node1593_l;
      node1595 = node1593_r;
      node1596_r = node1592_r & pixel[380];
      node1596_l = node1592_r & ~pixel[380];
      node1597 = node1596_l;
      node1598 = node1596_r;
      node1599_r = node1591_r & pixel[428];
      node1599_l = node1591_r & ~pixel[428];
      node1600_r = node1599_l & pixel[459];
      node1600_l = node1599_l & ~pixel[459];
      node1601 = node1600_l;
      node1602 = node1600_r;
      node1603_r = node1599_r & pixel[233];
      node1603_l = node1599_r & ~pixel[233];
      node1604 = node1603_l;
      node1605 = node1603_r;
      node1606_r = node1590_r & pixel[497];
      node1606_l = node1590_r & ~pixel[497];
      node1607 = node1606_l;
      node1608_r = node1606_r & pixel[155];
      node1608_l = node1606_r & ~pixel[155];
      node1609 = node1608_l;
      node1610_r = node1608_r & pixel[411];
      node1610_l = node1608_r & ~pixel[411];
      node1611 = node1610_l;
      node1612 = node1610_r;
      node1613_r = node1589_r & pixel[174];
      node1613_l = node1589_r & ~pixel[174];
      node1614_r = node1613_l & pixel[452];
      node1614_l = node1613_l & ~pixel[452];
      node1615_r = node1614_l & pixel[487];
      node1615_l = node1614_l & ~pixel[487];
      node1616_r = node1615_l & pixel[547];
      node1616_l = node1615_l & ~pixel[547];
      node1617 = node1616_l;
      node1618 = node1616_r;
      node1619_r = node1615_r & pixel[436];
      node1619_l = node1615_r & ~pixel[436];
      node1620 = node1619_l;
      node1621 = node1619_r;
      node1622 = node1614_r;
      node1623_r = node1613_r & pixel[485];
      node1623_l = node1613_r & ~pixel[485];
      node1624 = node1623_l;
      node1625_r = node1623_r & pixel[467];
      node1625_l = node1623_r & ~pixel[467];
      node1626 = node1625_l;
      node1627_r = node1625_r & pixel[258];
      node1627_l = node1625_r & ~pixel[258];
      node1628 = node1627_l;
      node1629 = node1627_r;
      node1630_r = node1524_r & pixel[460];
      node1630_l = node1524_r & ~pixel[460];
      node1631_r = node1630_l & pixel[357];
      node1631_l = node1630_l & ~pixel[357];
      node1632_r = node1631_l & pixel[429];
      node1632_l = node1631_l & ~pixel[429];
      node1633_r = node1632_l & pixel[459];
      node1633_l = node1632_l & ~pixel[459];
      node1634_r = node1633_l & pixel[439];
      node1634_l = node1633_l & ~pixel[439];
      node1635_r = node1634_l & pixel[345];
      node1635_l = node1634_l & ~pixel[345];
      node1636 = node1635_l;
      node1637 = node1635_r;
      node1638_r = node1634_r & pixel[666];
      node1638_l = node1634_r & ~pixel[666];
      node1639 = node1638_l;
      node1640 = node1638_r;
      node1641_r = node1633_r & pixel[147];
      node1641_l = node1633_r & ~pixel[147];
      node1642_r = node1641_l & pixel[245];
      node1642_l = node1641_l & ~pixel[245];
      node1643 = node1642_l;
      node1644 = node1642_r;
      node1645 = node1641_r;
      node1646_r = node1632_r & pixel[405];
      node1646_l = node1632_r & ~pixel[405];
      node1647_r = node1646_l & pixel[406];
      node1647_l = node1646_l & ~pixel[406];
      node1648_r = node1647_l & pixel[383];
      node1648_l = node1647_l & ~pixel[383];
      node1649 = node1648_l;
      node1650 = node1648_r;
      node1651_r = node1647_r & pixel[456];
      node1651_l = node1647_r & ~pixel[456];
      node1652 = node1651_l;
      node1653 = node1651_r;
      node1654_r = node1646_r & pixel[352];
      node1654_l = node1646_r & ~pixel[352];
      node1655_r = node1654_l & pixel[236];
      node1655_l = node1654_l & ~pixel[236];
      node1656 = node1655_l;
      node1657 = node1655_r;
      node1658_r = node1654_r & pixel[651];
      node1658_l = node1654_r & ~pixel[651];
      node1659 = node1658_l;
      node1660 = node1658_r;
      node1661_r = node1631_r & pixel[264];
      node1661_l = node1631_r & ~pixel[264];
      node1662_r = node1661_l & pixel[536];
      node1662_l = node1661_l & ~pixel[536];
      node1663_r = node1662_l & pixel[121];
      node1663_l = node1662_l & ~pixel[121];
      node1664_r = node1663_l & pixel[575];
      node1664_l = node1663_l & ~pixel[575];
      node1665 = node1664_l;
      node1666 = node1664_r;
      node1667_r = node1663_r & pixel[608];
      node1667_l = node1663_r & ~pixel[608];
      node1668 = node1667_l;
      node1669 = node1667_r;
      node1670 = node1662_r;
      node1671_r = node1661_r & pixel[429];
      node1671_l = node1661_r & ~pixel[429];
      node1672_r = node1671_l & pixel[426];
      node1672_l = node1671_l & ~pixel[426];
      node1673_r = node1672_l & pixel[653];
      node1673_l = node1672_l & ~pixel[653];
      node1674 = node1673_l;
      node1675 = node1673_r;
      node1676 = node1672_r;
      node1677_r = node1671_r & pixel[203];
      node1677_l = node1671_r & ~pixel[203];
      node1678_r = node1677_l & pixel[468];
      node1678_l = node1677_l & ~pixel[468];
      node1679 = node1678_l;
      node1680 = node1678_r;
      node1681_r = node1677_r & pixel[159];
      node1681_l = node1677_r & ~pixel[159];
      node1682 = node1681_l;
      node1683 = node1681_r;
      node1684_r = node1630_r & pixel[584];
      node1684_l = node1630_r & ~pixel[584];
      node1685_r = node1684_l & pixel[428];
      node1685_l = node1684_l & ~pixel[428];
      node1686_r = node1685_l & pixel[406];
      node1686_l = node1685_l & ~pixel[406];
      node1687_r = node1686_l & pixel[490];
      node1687_l = node1686_l & ~pixel[490];
      node1688_r = node1687_l & pixel[655];
      node1688_l = node1687_l & ~pixel[655];
      node1689 = node1688_l;
      node1690 = node1688_r;
      node1691_r = node1687_r & pixel[128];
      node1691_l = node1687_r & ~pixel[128];
      node1692 = node1691_l;
      node1693 = node1691_r;
      node1694_r = node1686_r & pixel[638];
      node1694_l = node1686_r & ~pixel[638];
      node1695_r = node1694_l & pixel[130];
      node1695_l = node1694_l & ~pixel[130];
      node1696 = node1695_l;
      node1697 = node1695_r;
      node1698_r = node1694_r & pixel[688];
      node1698_l = node1694_r & ~pixel[688];
      node1699 = node1698_l;
      node1700 = node1698_r;
      node1701_r = node1685_r & pixel[381];
      node1701_l = node1685_r & ~pixel[381];
      node1702_r = node1701_l & pixel[385];
      node1702_l = node1701_l & ~pixel[385];
      node1703_r = node1702_l & pixel[600];
      node1703_l = node1702_l & ~pixel[600];
      node1704 = node1703_l;
      node1705 = node1703_r;
      node1706_r = node1702_r & pixel[409];
      node1706_l = node1702_r & ~pixel[409];
      node1707 = node1706_l;
      node1708 = node1706_r;
      node1709_r = node1701_r & pixel[597];
      node1709_l = node1701_r & ~pixel[597];
      node1710_r = node1709_l & pixel[183];
      node1710_l = node1709_l & ~pixel[183];
      node1711 = node1710_l;
      node1712 = node1710_r;
      node1713_r = node1709_r & pixel[408];
      node1713_l = node1709_r & ~pixel[408];
      node1714 = node1713_l;
      node1715 = node1713_r;
      node1716_r = node1684_r & pixel[330];
      node1716_l = node1684_r & ~pixel[330];
      node1717_r = node1716_l & pixel[325];
      node1717_l = node1716_l & ~pixel[325];
      node1718 = node1717_l;
      node1719 = node1717_r;
      node1720_r = node1716_r & pixel[145];
      node1720_l = node1716_r & ~pixel[145];
      node1721 = node1720_l;
      node1722_r = node1720_r & pixel[285];
      node1722_l = node1720_r & ~pixel[285];
      node1723 = node1722_l;
      node1724 = node1722_r;
      result0 = node75 | node89 | node108 | node135 | node138 | node147 | node217 | node226 | node255 | node263 | node270 | node276 | node277 | node283 | node288 | node296 | node301 | node302 | node310 | node320 | node324 | node330 | node331 | node333 | node341 | node342 | node345 | node349 | node350 | node352 | node355 | node359 | node369 | node381 | node390 | node393 | node446 | node456 | node541 | node564 | node611 | node639 | node671 | node741 | node745 | node746 | node751 | node790 | node807 | node822 | node883 | node929 | node942 | node982 | node999 | node1011 | node1014 | node1022 | node1046 | node1051 | node1071 | node1086 | node1089 | node1090 | node1111 | node1112 | node1115 | node1136 | node1141 | node1151 | node1158 | node1160 | node1161 | node1165 | node1172 | node1173 | node1175 | node1187 | node1211 | node1222 | node1226 | node1227 | node1241 | node1261 | node1266 | node1281 | node1285 | node1289 | node1299 | node1301 | node1320 | node1321 | node1338 | node1343 | node1344 | node1346 | node1347 | node1354 | node1360 | node1362 | node1365 | node1371 | node1372 | node1376 | node1377 | node1380 | node1385 | node1387 | node1388 | node1395 | node1413 | node1416 | node1460 | node1472 | node1480 | node1494 | node1521 | node1609 | node1650 | node1656 | node1666 | node1676 | node1679 | node1680 | node1682 | node1690 | node1693 | node1707 | node1708 | node1714 | node1723;
      result1 = node10 | node25 | node48 | node170 | node259 | node409 | node804 | node812 | node873 | node888 | node889 | node891 | node898;
      result2 = node11 | node18 | node20 | node26 | node32 | node42 | node45 | node56 | node57 | node78 | node83 | node86 | node243 | node274 | node280 | node308 | node344 | node365 | node370 | node378 | node387 | node447 | node451 | node452 | node453 | node472 | node480 | node484 | node488 | node493 | node554 | node568 | node571 | node576 | node578 | node593 | node596 | node607 | node608 | node631 | node640 | node672 | node685 | node725 | node726 | node730 | node739 | node742 | node757 | node821 | node832 | node876 | node884 | node904 | node905 | node908 | node911 | node912 | node914 | node915 | node919 | node930 | node936 | node937 | node949 | node950 | node954 | node957 | node958 | node963 | node964 | node970 | node980 | node991 | node998 | node1003 | node1015 | node1018 | node1026 | node1027 | node1043 | node1044 | node1057 | node1064 | node1079 | node1102 | node1106 | node1178 | node1189 | node1202 | node1204 | node1232 | node1253 | node1262 | node1275 | node1276 | node1298 | node1302 | node1305 | node1309 | node1326 | node1327 | node1359 | node1373 | node1409 | node1423 | node1424 | node1427 | node1434 | node1438 | node1452 | node1453 | node1455 | node1458 | node1466 | node1469 | node1503 | node1510 | node1538 | node1541 | node1556 | node1565 | node1569 | node1587 | node1588 | node1669 | node1699 | node1719 | node1724;
      result3 = node13 | node35 | node41 | node44 | node51 | node77 | node90 | node92 | node120 | node134 | node139 | node141 | node173 | node177 | node256 | node260 | node273 | node287 | node293 | node294 | node305 | node307 | node373 | node408 | node437 | node439 | node440 | node444 | node487 | node535 | node553 | node556 | node557 | node561 | node603 | node648 | node651 | node652 | node703 | node710 | node729 | node732 | node755 | node775 | node784 | node787 | node796 | node806 | node811 | node814 | node818 | node819 | node829 | node831 | node843 | node850 | node853 | node854 | node858 | node945 | node951 | node955 | node1098 | node1168 | node1180 | node1235 | node1246 | node1247 | node1250 | node1257 | node1278 | node1296 | node1306 | node1311 | node1331 | node1350 | node1358 | node1364 | node1392 | node1456 | node1531 | node1539 | node1542 | node1547 | node1553 | node1554 | node1566 | node1570 | node1580 | node1584 | node1585 | node1598 | node1618 | node1624 | node1628 | node1636 | node1639 | node1645 | node1660 | node1668 | node1670 | node1674 | node1683 | node1689 | node1704;
      result4 = node106 | node163 | node241 | node244 | node247 | node323 | node367 | node386 | node392 | node406 | node416 | node420 | node424 | node431 | node463 | node465 | node466 | node473 | node511 | node512 | node544 | node585 | node600 | node616 | node617 | node619 | node624 | node677 | node709 | node716 | node738 | node748 | node768 | node772 | node781 | node797 | node799 | node800 | node803 | node828 | node836 | node839 | node861 | node863 | node966 | node994 | node1006 | node1034 | node1037 | node1053 | node1059 | node1067 | node1072 | node1075 | node1130 | node1134 | node1148 | node1201 | node1209 | node1236 | node1239 | node1439 | node1465 | node1486 | node1491 | node1507 | node1522 | node1711;
      result5 = node29 | node49 | node62 | node72 | node98 | node101 | node116 | node131 | node142 | node146 | node150 | node153 | node156 | node157 | node162 | node178 | node191 | node194 | node196 | node198 | node202 | node204 | node207 | node212 | node216 | node225 | node228 | node235 | node240 | node254 | node261 | node265 | node282 | node286 | node299 | node311 | node335 | node347 | node436 | node443 | node478 | node509 | node525 | node548 | node560 | node595 | node637 | node649 | node656 | node657 | node661 | node662 | node664 | node665 | node678 | node692 | node696 | node700 | node769 | node788 | node791 | node838 | node844 | node862 | node941 | node979 | node1002 | node1114 | node1128 | node1140 | node1143 | node1157 | node1164 | node1167 | node1176 | node1194 | node1220 | node1256 | node1280 | node1295 | node1332 | node1336 | node1337 | node1379 | node1384 | node1391 | node1394 | node1402 | node1404 | node1482 | node1499 | node1500 | node1515 | node1534 | node1535 | node1546 | node1549 | node1550 | node1557 | node1577 | node1594 | node1595 | node1597 | node1601 | node1605 | node1612 | node1622 | node1626 | node1637 | node1640 | node1657 | node1705 | node1718;
      result6 = node58 | node60 | node105 | node132 | node154 | node181 | node187 | node377 | node384 | node412 | node430 | node455 | node462 | node477 | node636 | node680 | node681 | node684 | node874 | node877 | node880 | node881 | node920 | node922 | node926 | node927 | node944 | node967 | node976 | node983 | node990 | node993 | node997 | node1021 | node1033 | node1054 | node1074 | node1099 | node1101 | node1105 | node1107 | node1118 | node1119 | node1181 | node1208 | node1212 | node1219 | node1223 | node1228 | node1233 | node1240 | node1249 | node1254 | node1263 | node1267 | node1268 | node1273 | node1284 | node1287 | node1290 | node1310 | node1322 | node1353 | node1461 | node1478 | node1563 | node1578 | node1604 | node1611 | node1652;
      result7 = node17 | node33 | node69 | node70 | node73 | node82 | node93 | node102 | node113 | node149 | node229 | node232 | node318 | node329 | node405 | node413 | node423 | node427 | node469 | node496 | node501 | node503 | node515 | node517 | node524 | node527 | node528 | node532 | node534 | node540 | node620 | node627 | node633 | node688 | node765 | node835 | node846 | node859 | node895 | node938 | node1012 | node1065 | node1082 | node1135 | node1150 | node1190 | node1196 | node1426 | node1430 | node1431 | node1441 | node1446;
      result8 = node14 | node28 | node36 | node52 | node63 | node85 | node109 | node117 | node123 | node166 | node169 | node172 | node180 | node184 | node185 | node188 | node197 | node205 | node208 | node213 | node215 | node248 | node266 | node297 | node336 | node356 | node358 | node366 | node380 | node395 | node428 | node481 | node485 | node569 | node572 | node575 | node579 | node669 | node687 | node693 | node695 | node699 | node702 | node717 | node719 | node733 | node749 | node754 | node758 | node776 | node783 | node815 | node847 | node851 | node892 | node896 | node899 | node907 | node923 | node974 | node1030 | node1122 | node1127 | node1131 | node1144 | node1147 | node1186 | node1193 | node1197 | node1205 | node1325 | node1333 | node1351 | node1400 | node1405 | node1410 | node1412 | node1415 | node1433 | node1447 | node1471 | node1479 | node1483 | node1487 | node1493 | node1502 | node1506 | node1509 | node1514 | node1517 | node1518 | node1532 | node1562 | node1572 | node1573 | node1581 | node1602 | node1607 | node1617 | node1620 | node1621 | node1629 | node1643 | node1644 | node1649 | node1653 | node1659 | node1665 | node1675 | node1692 | node1696 | node1697 | node1700 | node1712 | node1715 | node1721;
      result9 = node21 | node99 | node114 | node121 | node124 | node165 | node233 | node236 | node249 | node319 | node325 | node374 | node396 | node415 | node421 | node470 | node494 | node497 | node500 | node504 | node508 | node516 | node531 | node539 | node545 | node547 | node563 | node586 | node588 | node589 | node592 | node601 | node604 | node610 | node623 | node626 | node632 | node655 | node668 | node712 | node713 | node720 | node724 | node766 | node773 | node780 | node971 | node973 | node1005 | node1019 | node1029 | node1036 | node1047 | node1050 | node1058 | node1068 | node1080 | node1083 | node1087 | node1121 | node1401 | node1442 | node1445 | node1467 | node1490 | node1523;

      tree_7 = {result9, result8, result7, result6, result5, result4, result3, result2, result1, result0};
    end
  endfunction

  function [9:0] tree_8;
    input [783:0] pixel;

    reg node0_r;
    reg node0_l;
    reg node1_r;
    reg node1_l;
    reg node2_r;
    reg node2_l;
    reg node3_r;
    reg node3_l;
    reg node4_r;
    reg node4_l;
    reg node5_r;
    reg node5_l;
    reg node6_r;
    reg node6_l;
    reg node7_r;
    reg node7_l;
    reg node8_r;
    reg node8_l;
    reg node9_r;
    reg node9_l;
    reg node10;
    reg node11;
    reg node12_r;
    reg node12_l;
    reg node13;
    reg node14;
    reg node15_r;
    reg node15_l;
    reg node16_r;
    reg node16_l;
    reg node17;
    reg node18;
    reg node19_r;
    reg node19_l;
    reg node20;
    reg node21;
    reg node22_r;
    reg node22_l;
    reg node23_r;
    reg node23_l;
    reg node24_r;
    reg node24_l;
    reg node25;
    reg node26;
    reg node27_r;
    reg node27_l;
    reg node28;
    reg node29;
    reg node30_r;
    reg node30_l;
    reg node31_r;
    reg node31_l;
    reg node32;
    reg node33;
    reg node34_r;
    reg node34_l;
    reg node35;
    reg node36;
    reg node37_r;
    reg node37_l;
    reg node38_r;
    reg node38_l;
    reg node39_r;
    reg node39_l;
    reg node40_r;
    reg node40_l;
    reg node41;
    reg node42;
    reg node43_r;
    reg node43_l;
    reg node44;
    reg node45;
    reg node46_r;
    reg node46_l;
    reg node47_r;
    reg node47_l;
    reg node48;
    reg node49;
    reg node50_r;
    reg node50_l;
    reg node51;
    reg node52;
    reg node53_r;
    reg node53_l;
    reg node54_r;
    reg node54_l;
    reg node55_r;
    reg node55_l;
    reg node56;
    reg node57;
    reg node58_r;
    reg node58_l;
    reg node59;
    reg node60;
    reg node61_r;
    reg node61_l;
    reg node62_r;
    reg node62_l;
    reg node63;
    reg node64;
    reg node65_r;
    reg node65_l;
    reg node66;
    reg node67;
    reg node68_r;
    reg node68_l;
    reg node69_r;
    reg node69_l;
    reg node70_r;
    reg node70_l;
    reg node71_r;
    reg node71_l;
    reg node72_r;
    reg node72_l;
    reg node73;
    reg node74;
    reg node75_r;
    reg node75_l;
    reg node76;
    reg node77;
    reg node78_r;
    reg node78_l;
    reg node79_r;
    reg node79_l;
    reg node80;
    reg node81;
    reg node82_r;
    reg node82_l;
    reg node83;
    reg node84;
    reg node85_r;
    reg node85_l;
    reg node86_r;
    reg node86_l;
    reg node87_r;
    reg node87_l;
    reg node88;
    reg node89;
    reg node90_r;
    reg node90_l;
    reg node91;
    reg node92;
    reg node93_r;
    reg node93_l;
    reg node94_r;
    reg node94_l;
    reg node95;
    reg node96;
    reg node97;
    reg node98_r;
    reg node98_l;
    reg node99_r;
    reg node99_l;
    reg node100_r;
    reg node100_l;
    reg node101_r;
    reg node101_l;
    reg node102;
    reg node103;
    reg node104;
    reg node105;
    reg node106_r;
    reg node106_l;
    reg node107_r;
    reg node107_l;
    reg node108_r;
    reg node108_l;
    reg node109;
    reg node110;
    reg node111_r;
    reg node111_l;
    reg node112;
    reg node113;
    reg node114;
    reg node115_r;
    reg node115_l;
    reg node116_r;
    reg node116_l;
    reg node117_r;
    reg node117_l;
    reg node118_r;
    reg node118_l;
    reg node119_r;
    reg node119_l;
    reg node120_r;
    reg node120_l;
    reg node121;
    reg node122;
    reg node123_r;
    reg node123_l;
    reg node124;
    reg node125;
    reg node126_r;
    reg node126_l;
    reg node127_r;
    reg node127_l;
    reg node128;
    reg node129;
    reg node130_r;
    reg node130_l;
    reg node131;
    reg node132;
    reg node133_r;
    reg node133_l;
    reg node134_r;
    reg node134_l;
    reg node135_r;
    reg node135_l;
    reg node136;
    reg node137;
    reg node138_r;
    reg node138_l;
    reg node139;
    reg node140;
    reg node141_r;
    reg node141_l;
    reg node142_r;
    reg node142_l;
    reg node143;
    reg node144;
    reg node145_r;
    reg node145_l;
    reg node146;
    reg node147;
    reg node148;
    reg node149_r;
    reg node149_l;
    reg node150_r;
    reg node150_l;
    reg node151_r;
    reg node151_l;
    reg node152_r;
    reg node152_l;
    reg node153_r;
    reg node153_l;
    reg node154;
    reg node155;
    reg node156_r;
    reg node156_l;
    reg node157;
    reg node158;
    reg node159_r;
    reg node159_l;
    reg node160_r;
    reg node160_l;
    reg node161;
    reg node162;
    reg node163_r;
    reg node163_l;
    reg node164;
    reg node165;
    reg node166_r;
    reg node166_l;
    reg node167_r;
    reg node167_l;
    reg node168_r;
    reg node168_l;
    reg node169;
    reg node170;
    reg node171_r;
    reg node171_l;
    reg node172;
    reg node173;
    reg node174_r;
    reg node174_l;
    reg node175_r;
    reg node175_l;
    reg node176;
    reg node177;
    reg node178_r;
    reg node178_l;
    reg node179;
    reg node180;
    reg node181_r;
    reg node181_l;
    reg node182_r;
    reg node182_l;
    reg node183_r;
    reg node183_l;
    reg node184_r;
    reg node184_l;
    reg node185;
    reg node186;
    reg node187_r;
    reg node187_l;
    reg node188;
    reg node189;
    reg node190_r;
    reg node190_l;
    reg node191_r;
    reg node191_l;
    reg node192;
    reg node193;
    reg node194;
    reg node195_r;
    reg node195_l;
    reg node196_r;
    reg node196_l;
    reg node197_r;
    reg node197_l;
    reg node198;
    reg node199;
    reg node200_r;
    reg node200_l;
    reg node201;
    reg node202;
    reg node203_r;
    reg node203_l;
    reg node204_r;
    reg node204_l;
    reg node205;
    reg node206;
    reg node207_r;
    reg node207_l;
    reg node208;
    reg node209;
    reg node210_r;
    reg node210_l;
    reg node211_r;
    reg node211_l;
    reg node212_r;
    reg node212_l;
    reg node213_r;
    reg node213_l;
    reg node214_r;
    reg node214_l;
    reg node215_r;
    reg node215_l;
    reg node216_r;
    reg node216_l;
    reg node217;
    reg node218;
    reg node219_r;
    reg node219_l;
    reg node220;
    reg node221;
    reg node222_r;
    reg node222_l;
    reg node223_r;
    reg node223_l;
    reg node224;
    reg node225;
    reg node226_r;
    reg node226_l;
    reg node227;
    reg node228;
    reg node229_r;
    reg node229_l;
    reg node230_r;
    reg node230_l;
    reg node231_r;
    reg node231_l;
    reg node232;
    reg node233;
    reg node234_r;
    reg node234_l;
    reg node235;
    reg node236;
    reg node237_r;
    reg node237_l;
    reg node238_r;
    reg node238_l;
    reg node239;
    reg node240;
    reg node241;
    reg node242_r;
    reg node242_l;
    reg node243_r;
    reg node243_l;
    reg node244_r;
    reg node244_l;
    reg node245_r;
    reg node245_l;
    reg node246;
    reg node247;
    reg node248_r;
    reg node248_l;
    reg node249;
    reg node250;
    reg node251_r;
    reg node251_l;
    reg node252_r;
    reg node252_l;
    reg node253;
    reg node254;
    reg node255;
    reg node256_r;
    reg node256_l;
    reg node257_r;
    reg node257_l;
    reg node258_r;
    reg node258_l;
    reg node259;
    reg node260;
    reg node261_r;
    reg node261_l;
    reg node262;
    reg node263;
    reg node264_r;
    reg node264_l;
    reg node265_r;
    reg node265_l;
    reg node266;
    reg node267;
    reg node268_r;
    reg node268_l;
    reg node269;
    reg node270;
    reg node271_r;
    reg node271_l;
    reg node272_r;
    reg node272_l;
    reg node273_r;
    reg node273_l;
    reg node274_r;
    reg node274_l;
    reg node275_r;
    reg node275_l;
    reg node276;
    reg node277;
    reg node278_r;
    reg node278_l;
    reg node279;
    reg node280;
    reg node281_r;
    reg node281_l;
    reg node282_r;
    reg node282_l;
    reg node283;
    reg node284;
    reg node285_r;
    reg node285_l;
    reg node286;
    reg node287;
    reg node288_r;
    reg node288_l;
    reg node289_r;
    reg node289_l;
    reg node290_r;
    reg node290_l;
    reg node291;
    reg node292;
    reg node293_r;
    reg node293_l;
    reg node294;
    reg node295;
    reg node296_r;
    reg node296_l;
    reg node297_r;
    reg node297_l;
    reg node298;
    reg node299;
    reg node300_r;
    reg node300_l;
    reg node301;
    reg node302;
    reg node303_r;
    reg node303_l;
    reg node304_r;
    reg node304_l;
    reg node305_r;
    reg node305_l;
    reg node306_r;
    reg node306_l;
    reg node307;
    reg node308;
    reg node309_r;
    reg node309_l;
    reg node310;
    reg node311;
    reg node312_r;
    reg node312_l;
    reg node313;
    reg node314;
    reg node315_r;
    reg node315_l;
    reg node316_r;
    reg node316_l;
    reg node317_r;
    reg node317_l;
    reg node318;
    reg node319;
    reg node320_r;
    reg node320_l;
    reg node321;
    reg node322;
    reg node323_r;
    reg node323_l;
    reg node324;
    reg node325_r;
    reg node325_l;
    reg node326;
    reg node327;
    reg node328_r;
    reg node328_l;
    reg node329_r;
    reg node329_l;
    reg node330_r;
    reg node330_l;
    reg node331_r;
    reg node331_l;
    reg node332_r;
    reg node332_l;
    reg node333_r;
    reg node333_l;
    reg node334;
    reg node335;
    reg node336_r;
    reg node336_l;
    reg node337;
    reg node338;
    reg node339_r;
    reg node339_l;
    reg node340_r;
    reg node340_l;
    reg node341;
    reg node342;
    reg node343_r;
    reg node343_l;
    reg node344;
    reg node345;
    reg node346_r;
    reg node346_l;
    reg node347_r;
    reg node347_l;
    reg node348_r;
    reg node348_l;
    reg node349;
    reg node350;
    reg node351_r;
    reg node351_l;
    reg node352;
    reg node353;
    reg node354_r;
    reg node354_l;
    reg node355_r;
    reg node355_l;
    reg node356;
    reg node357;
    reg node358_r;
    reg node358_l;
    reg node359;
    reg node360;
    reg node361_r;
    reg node361_l;
    reg node362_r;
    reg node362_l;
    reg node363_r;
    reg node363_l;
    reg node364_r;
    reg node364_l;
    reg node365;
    reg node366;
    reg node367_r;
    reg node367_l;
    reg node368;
    reg node369;
    reg node370_r;
    reg node370_l;
    reg node371_r;
    reg node371_l;
    reg node372;
    reg node373;
    reg node374;
    reg node375_r;
    reg node375_l;
    reg node376_r;
    reg node376_l;
    reg node377_r;
    reg node377_l;
    reg node378;
    reg node379;
    reg node380;
    reg node381;
    reg node382_r;
    reg node382_l;
    reg node383_r;
    reg node383_l;
    reg node384_r;
    reg node384_l;
    reg node385_r;
    reg node385_l;
    reg node386_r;
    reg node386_l;
    reg node387;
    reg node388;
    reg node389_r;
    reg node389_l;
    reg node390;
    reg node391;
    reg node392;
    reg node393_r;
    reg node393_l;
    reg node394_r;
    reg node394_l;
    reg node395_r;
    reg node395_l;
    reg node396;
    reg node397;
    reg node398_r;
    reg node398_l;
    reg node399;
    reg node400;
    reg node401_r;
    reg node401_l;
    reg node402;
    reg node403_r;
    reg node403_l;
    reg node404;
    reg node405;
    reg node406_r;
    reg node406_l;
    reg node407;
    reg node408;
    reg node409_r;
    reg node409_l;
    reg node410_r;
    reg node410_l;
    reg node411_r;
    reg node411_l;
    reg node412_r;
    reg node412_l;
    reg node413_r;
    reg node413_l;
    reg node414_r;
    reg node414_l;
    reg node415_r;
    reg node415_l;
    reg node416_r;
    reg node416_l;
    reg node417;
    reg node418;
    reg node419_r;
    reg node419_l;
    reg node420;
    reg node421;
    reg node422_r;
    reg node422_l;
    reg node423_r;
    reg node423_l;
    reg node424;
    reg node425;
    reg node426_r;
    reg node426_l;
    reg node427;
    reg node428;
    reg node429_r;
    reg node429_l;
    reg node430_r;
    reg node430_l;
    reg node431_r;
    reg node431_l;
    reg node432;
    reg node433;
    reg node434_r;
    reg node434_l;
    reg node435;
    reg node436;
    reg node437_r;
    reg node437_l;
    reg node438_r;
    reg node438_l;
    reg node439;
    reg node440;
    reg node441_r;
    reg node441_l;
    reg node442;
    reg node443;
    reg node444_r;
    reg node444_l;
    reg node445_r;
    reg node445_l;
    reg node446_r;
    reg node446_l;
    reg node447_r;
    reg node447_l;
    reg node448;
    reg node449;
    reg node450_r;
    reg node450_l;
    reg node451;
    reg node452;
    reg node453_r;
    reg node453_l;
    reg node454_r;
    reg node454_l;
    reg node455;
    reg node456;
    reg node457_r;
    reg node457_l;
    reg node458;
    reg node459;
    reg node460_r;
    reg node460_l;
    reg node461_r;
    reg node461_l;
    reg node462_r;
    reg node462_l;
    reg node463;
    reg node464;
    reg node465;
    reg node466_r;
    reg node466_l;
    reg node467;
    reg node468_r;
    reg node468_l;
    reg node469;
    reg node470;
    reg node471_r;
    reg node471_l;
    reg node472_r;
    reg node472_l;
    reg node473_r;
    reg node473_l;
    reg node474_r;
    reg node474_l;
    reg node475_r;
    reg node475_l;
    reg node476;
    reg node477;
    reg node478_r;
    reg node478_l;
    reg node479;
    reg node480;
    reg node481_r;
    reg node481_l;
    reg node482_r;
    reg node482_l;
    reg node483;
    reg node484;
    reg node485_r;
    reg node485_l;
    reg node486;
    reg node487;
    reg node488_r;
    reg node488_l;
    reg node489_r;
    reg node489_l;
    reg node490_r;
    reg node490_l;
    reg node491;
    reg node492;
    reg node493_r;
    reg node493_l;
    reg node494;
    reg node495;
    reg node496_r;
    reg node496_l;
    reg node497_r;
    reg node497_l;
    reg node498;
    reg node499;
    reg node500;
    reg node501_r;
    reg node501_l;
    reg node502_r;
    reg node502_l;
    reg node503_r;
    reg node503_l;
    reg node504_r;
    reg node504_l;
    reg node505;
    reg node506;
    reg node507_r;
    reg node507_l;
    reg node508;
    reg node509;
    reg node510_r;
    reg node510_l;
    reg node511_r;
    reg node511_l;
    reg node512;
    reg node513;
    reg node514_r;
    reg node514_l;
    reg node515;
    reg node516;
    reg node517_r;
    reg node517_l;
    reg node518_r;
    reg node518_l;
    reg node519_r;
    reg node519_l;
    reg node520;
    reg node521;
    reg node522_r;
    reg node522_l;
    reg node523;
    reg node524;
    reg node525_r;
    reg node525_l;
    reg node526_r;
    reg node526_l;
    reg node527;
    reg node528;
    reg node529_r;
    reg node529_l;
    reg node530;
    reg node531;
    reg node532_r;
    reg node532_l;
    reg node533_r;
    reg node533_l;
    reg node534_r;
    reg node534_l;
    reg node535_r;
    reg node535_l;
    reg node536_r;
    reg node536_l;
    reg node537_r;
    reg node537_l;
    reg node538;
    reg node539;
    reg node540_r;
    reg node540_l;
    reg node541;
    reg node542;
    reg node543_r;
    reg node543_l;
    reg node544;
    reg node545_r;
    reg node545_l;
    reg node546;
    reg node547;
    reg node548_r;
    reg node548_l;
    reg node549_r;
    reg node549_l;
    reg node550_r;
    reg node550_l;
    reg node551;
    reg node552;
    reg node553_r;
    reg node553_l;
    reg node554;
    reg node555;
    reg node556_r;
    reg node556_l;
    reg node557_r;
    reg node557_l;
    reg node558;
    reg node559;
    reg node560;
    reg node561_r;
    reg node561_l;
    reg node562_r;
    reg node562_l;
    reg node563_r;
    reg node563_l;
    reg node564_r;
    reg node564_l;
    reg node565;
    reg node566;
    reg node567_r;
    reg node567_l;
    reg node568;
    reg node569;
    reg node570_r;
    reg node570_l;
    reg node571_r;
    reg node571_l;
    reg node572;
    reg node573;
    reg node574;
    reg node575_r;
    reg node575_l;
    reg node576_r;
    reg node576_l;
    reg node577_r;
    reg node577_l;
    reg node578;
    reg node579;
    reg node580_r;
    reg node580_l;
    reg node581;
    reg node582;
    reg node583_r;
    reg node583_l;
    reg node584_r;
    reg node584_l;
    reg node585;
    reg node586;
    reg node587_r;
    reg node587_l;
    reg node588;
    reg node589;
    reg node590_r;
    reg node590_l;
    reg node591_r;
    reg node591_l;
    reg node592_r;
    reg node592_l;
    reg node593_r;
    reg node593_l;
    reg node594_r;
    reg node594_l;
    reg node595;
    reg node596;
    reg node597;
    reg node598_r;
    reg node598_l;
    reg node599_r;
    reg node599_l;
    reg node600;
    reg node601;
    reg node602;
    reg node603_r;
    reg node603_l;
    reg node604_r;
    reg node604_l;
    reg node605_r;
    reg node605_l;
    reg node606;
    reg node607;
    reg node608_r;
    reg node608_l;
    reg node609;
    reg node610;
    reg node611_r;
    reg node611_l;
    reg node612_r;
    reg node612_l;
    reg node613;
    reg node614;
    reg node615_r;
    reg node615_l;
    reg node616;
    reg node617;
    reg node618_r;
    reg node618_l;
    reg node619_r;
    reg node619_l;
    reg node620_r;
    reg node620_l;
    reg node621_r;
    reg node621_l;
    reg node622;
    reg node623;
    reg node624_r;
    reg node624_l;
    reg node625;
    reg node626;
    reg node627;
    reg node628_r;
    reg node628_l;
    reg node629_r;
    reg node629_l;
    reg node630;
    reg node631;
    reg node632_r;
    reg node632_l;
    reg node633_r;
    reg node633_l;
    reg node634;
    reg node635;
    reg node636;
    reg node637_r;
    reg node637_l;
    reg node638_r;
    reg node638_l;
    reg node639_r;
    reg node639_l;
    reg node640_r;
    reg node640_l;
    reg node641_r;
    reg node641_l;
    reg node642_r;
    reg node642_l;
    reg node643_r;
    reg node643_l;
    reg node644;
    reg node645;
    reg node646_r;
    reg node646_l;
    reg node647;
    reg node648;
    reg node649_r;
    reg node649_l;
    reg node650_r;
    reg node650_l;
    reg node651;
    reg node652;
    reg node653_r;
    reg node653_l;
    reg node654;
    reg node655;
    reg node656_r;
    reg node656_l;
    reg node657_r;
    reg node657_l;
    reg node658;
    reg node659_r;
    reg node659_l;
    reg node660;
    reg node661;
    reg node662_r;
    reg node662_l;
    reg node663_r;
    reg node663_l;
    reg node664;
    reg node665;
    reg node666;
    reg node667_r;
    reg node667_l;
    reg node668_r;
    reg node668_l;
    reg node669_r;
    reg node669_l;
    reg node670_r;
    reg node670_l;
    reg node671;
    reg node672;
    reg node673_r;
    reg node673_l;
    reg node674;
    reg node675;
    reg node676_r;
    reg node676_l;
    reg node677_r;
    reg node677_l;
    reg node678;
    reg node679;
    reg node680_r;
    reg node680_l;
    reg node681;
    reg node682;
    reg node683_r;
    reg node683_l;
    reg node684_r;
    reg node684_l;
    reg node685_r;
    reg node685_l;
    reg node686;
    reg node687;
    reg node688_r;
    reg node688_l;
    reg node689;
    reg node690;
    reg node691_r;
    reg node691_l;
    reg node692;
    reg node693;
    reg node694_r;
    reg node694_l;
    reg node695_r;
    reg node695_l;
    reg node696_r;
    reg node696_l;
    reg node697_r;
    reg node697_l;
    reg node698_r;
    reg node698_l;
    reg node699;
    reg node700;
    reg node701_r;
    reg node701_l;
    reg node702;
    reg node703;
    reg node704_r;
    reg node704_l;
    reg node705_r;
    reg node705_l;
    reg node706;
    reg node707;
    reg node708_r;
    reg node708_l;
    reg node709;
    reg node710;
    reg node711_r;
    reg node711_l;
    reg node712_r;
    reg node712_l;
    reg node713_r;
    reg node713_l;
    reg node714;
    reg node715;
    reg node716_r;
    reg node716_l;
    reg node717;
    reg node718;
    reg node719_r;
    reg node719_l;
    reg node720;
    reg node721;
    reg node722_r;
    reg node722_l;
    reg node723_r;
    reg node723_l;
    reg node724_r;
    reg node724_l;
    reg node725_r;
    reg node725_l;
    reg node726;
    reg node727;
    reg node728;
    reg node729_r;
    reg node729_l;
    reg node730_r;
    reg node730_l;
    reg node731;
    reg node732;
    reg node733_r;
    reg node733_l;
    reg node734;
    reg node735;
    reg node736_r;
    reg node736_l;
    reg node737_r;
    reg node737_l;
    reg node738_r;
    reg node738_l;
    reg node739;
    reg node740;
    reg node741_r;
    reg node741_l;
    reg node742;
    reg node743;
    reg node744_r;
    reg node744_l;
    reg node745_r;
    reg node745_l;
    reg node746;
    reg node747;
    reg node748_r;
    reg node748_l;
    reg node749;
    reg node750;
    reg node751_r;
    reg node751_l;
    reg node752_r;
    reg node752_l;
    reg node753_r;
    reg node753_l;
    reg node754_r;
    reg node754_l;
    reg node755_r;
    reg node755_l;
    reg node756_r;
    reg node756_l;
    reg node757;
    reg node758;
    reg node759_r;
    reg node759_l;
    reg node760;
    reg node761;
    reg node762_r;
    reg node762_l;
    reg node763_r;
    reg node763_l;
    reg node764;
    reg node765;
    reg node766_r;
    reg node766_l;
    reg node767;
    reg node768;
    reg node769_r;
    reg node769_l;
    reg node770;
    reg node771_r;
    reg node771_l;
    reg node772;
    reg node773_r;
    reg node773_l;
    reg node774;
    reg node775;
    reg node776_r;
    reg node776_l;
    reg node777_r;
    reg node777_l;
    reg node778_r;
    reg node778_l;
    reg node779_r;
    reg node779_l;
    reg node780;
    reg node781;
    reg node782_r;
    reg node782_l;
    reg node783;
    reg node784;
    reg node785_r;
    reg node785_l;
    reg node786_r;
    reg node786_l;
    reg node787;
    reg node788;
    reg node789;
    reg node790_r;
    reg node790_l;
    reg node791_r;
    reg node791_l;
    reg node792_r;
    reg node792_l;
    reg node793;
    reg node794;
    reg node795_r;
    reg node795_l;
    reg node796;
    reg node797;
    reg node798_r;
    reg node798_l;
    reg node799_r;
    reg node799_l;
    reg node800;
    reg node801;
    reg node802_r;
    reg node802_l;
    reg node803;
    reg node804;
    reg node805_r;
    reg node805_l;
    reg node806_r;
    reg node806_l;
    reg node807_r;
    reg node807_l;
    reg node808_r;
    reg node808_l;
    reg node809_r;
    reg node809_l;
    reg node810;
    reg node811;
    reg node812_r;
    reg node812_l;
    reg node813;
    reg node814;
    reg node815_r;
    reg node815_l;
    reg node816_r;
    reg node816_l;
    reg node817;
    reg node818;
    reg node819_r;
    reg node819_l;
    reg node820;
    reg node821;
    reg node822_r;
    reg node822_l;
    reg node823_r;
    reg node823_l;
    reg node824_r;
    reg node824_l;
    reg node825;
    reg node826;
    reg node827_r;
    reg node827_l;
    reg node828;
    reg node829;
    reg node830_r;
    reg node830_l;
    reg node831_r;
    reg node831_l;
    reg node832;
    reg node833;
    reg node834_r;
    reg node834_l;
    reg node835;
    reg node836;
    reg node837_r;
    reg node837_l;
    reg node838_r;
    reg node838_l;
    reg node839_r;
    reg node839_l;
    reg node840_r;
    reg node840_l;
    reg node841;
    reg node842;
    reg node843_r;
    reg node843_l;
    reg node844;
    reg node845;
    reg node846_r;
    reg node846_l;
    reg node847_r;
    reg node847_l;
    reg node848;
    reg node849;
    reg node850_r;
    reg node850_l;
    reg node851;
    reg node852;
    reg node853_r;
    reg node853_l;
    reg node854_r;
    reg node854_l;
    reg node855_r;
    reg node855_l;
    reg node856;
    reg node857;
    reg node858_r;
    reg node858_l;
    reg node859;
    reg node860;
    reg node861_r;
    reg node861_l;
    reg node862_r;
    reg node862_l;
    reg node863;
    reg node864;
    reg node865;
    reg node866_r;
    reg node866_l;
    reg node867_r;
    reg node867_l;
    reg node868_r;
    reg node868_l;
    reg node869_r;
    reg node869_l;
    reg node870_r;
    reg node870_l;
    reg node871_r;
    reg node871_l;
    reg node872_r;
    reg node872_l;
    reg node873_r;
    reg node873_l;
    reg node874_r;
    reg node874_l;
    reg node875;
    reg node876;
    reg node877_r;
    reg node877_l;
    reg node878;
    reg node879;
    reg node880_r;
    reg node880_l;
    reg node881_r;
    reg node881_l;
    reg node882;
    reg node883;
    reg node884_r;
    reg node884_l;
    reg node885;
    reg node886;
    reg node887_r;
    reg node887_l;
    reg node888_r;
    reg node888_l;
    reg node889_r;
    reg node889_l;
    reg node890;
    reg node891;
    reg node892_r;
    reg node892_l;
    reg node893;
    reg node894;
    reg node895_r;
    reg node895_l;
    reg node896_r;
    reg node896_l;
    reg node897;
    reg node898;
    reg node899_r;
    reg node899_l;
    reg node900;
    reg node901;
    reg node902_r;
    reg node902_l;
    reg node903_r;
    reg node903_l;
    reg node904_r;
    reg node904_l;
    reg node905_r;
    reg node905_l;
    reg node906;
    reg node907;
    reg node908_r;
    reg node908_l;
    reg node909;
    reg node910;
    reg node911_r;
    reg node911_l;
    reg node912_r;
    reg node912_l;
    reg node913;
    reg node914;
    reg node915_r;
    reg node915_l;
    reg node916;
    reg node917;
    reg node918_r;
    reg node918_l;
    reg node919_r;
    reg node919_l;
    reg node920_r;
    reg node920_l;
    reg node921;
    reg node922;
    reg node923_r;
    reg node923_l;
    reg node924;
    reg node925;
    reg node926_r;
    reg node926_l;
    reg node927_r;
    reg node927_l;
    reg node928;
    reg node929;
    reg node930;
    reg node931_r;
    reg node931_l;
    reg node932_r;
    reg node932_l;
    reg node933_r;
    reg node933_l;
    reg node934_r;
    reg node934_l;
    reg node935_r;
    reg node935_l;
    reg node936;
    reg node937;
    reg node938_r;
    reg node938_l;
    reg node939;
    reg node940;
    reg node941_r;
    reg node941_l;
    reg node942_r;
    reg node942_l;
    reg node943;
    reg node944;
    reg node945_r;
    reg node945_l;
    reg node946;
    reg node947;
    reg node948_r;
    reg node948_l;
    reg node949_r;
    reg node949_l;
    reg node950_r;
    reg node950_l;
    reg node951;
    reg node952;
    reg node953_r;
    reg node953_l;
    reg node954;
    reg node955;
    reg node956_r;
    reg node956_l;
    reg node957_r;
    reg node957_l;
    reg node958;
    reg node959;
    reg node960_r;
    reg node960_l;
    reg node961;
    reg node962;
    reg node963_r;
    reg node963_l;
    reg node964_r;
    reg node964_l;
    reg node965_r;
    reg node965_l;
    reg node966_r;
    reg node966_l;
    reg node967;
    reg node968;
    reg node969_r;
    reg node969_l;
    reg node970;
    reg node971;
    reg node972_r;
    reg node972_l;
    reg node973_r;
    reg node973_l;
    reg node974;
    reg node975;
    reg node976_r;
    reg node976_l;
    reg node977;
    reg node978;
    reg node979_r;
    reg node979_l;
    reg node980_r;
    reg node980_l;
    reg node981_r;
    reg node981_l;
    reg node982;
    reg node983;
    reg node984_r;
    reg node984_l;
    reg node985;
    reg node986;
    reg node987_r;
    reg node987_l;
    reg node988_r;
    reg node988_l;
    reg node989;
    reg node990;
    reg node991_r;
    reg node991_l;
    reg node992;
    reg node993;
    reg node994_r;
    reg node994_l;
    reg node995_r;
    reg node995_l;
    reg node996_r;
    reg node996_l;
    reg node997_r;
    reg node997_l;
    reg node998_r;
    reg node998_l;
    reg node999_r;
    reg node999_l;
    reg node1000;
    reg node1001;
    reg node1002_r;
    reg node1002_l;
    reg node1003;
    reg node1004;
    reg node1005_r;
    reg node1005_l;
    reg node1006_r;
    reg node1006_l;
    reg node1007;
    reg node1008;
    reg node1009_r;
    reg node1009_l;
    reg node1010;
    reg node1011;
    reg node1012_r;
    reg node1012_l;
    reg node1013_r;
    reg node1013_l;
    reg node1014_r;
    reg node1014_l;
    reg node1015;
    reg node1016;
    reg node1017_r;
    reg node1017_l;
    reg node1018;
    reg node1019;
    reg node1020_r;
    reg node1020_l;
    reg node1021;
    reg node1022_r;
    reg node1022_l;
    reg node1023;
    reg node1024;
    reg node1025_r;
    reg node1025_l;
    reg node1026_r;
    reg node1026_l;
    reg node1027_r;
    reg node1027_l;
    reg node1028_r;
    reg node1028_l;
    reg node1029;
    reg node1030;
    reg node1031_r;
    reg node1031_l;
    reg node1032;
    reg node1033;
    reg node1034_r;
    reg node1034_l;
    reg node1035;
    reg node1036_r;
    reg node1036_l;
    reg node1037;
    reg node1038;
    reg node1039_r;
    reg node1039_l;
    reg node1040_r;
    reg node1040_l;
    reg node1041_r;
    reg node1041_l;
    reg node1042;
    reg node1043;
    reg node1044;
    reg node1045_r;
    reg node1045_l;
    reg node1046_r;
    reg node1046_l;
    reg node1047;
    reg node1048;
    reg node1049_r;
    reg node1049_l;
    reg node1050;
    reg node1051;
    reg node1052_r;
    reg node1052_l;
    reg node1053_r;
    reg node1053_l;
    reg node1054_r;
    reg node1054_l;
    reg node1055_r;
    reg node1055_l;
    reg node1056_r;
    reg node1056_l;
    reg node1057;
    reg node1058;
    reg node1059_r;
    reg node1059_l;
    reg node1060;
    reg node1061;
    reg node1062_r;
    reg node1062_l;
    reg node1063_r;
    reg node1063_l;
    reg node1064;
    reg node1065;
    reg node1066_r;
    reg node1066_l;
    reg node1067;
    reg node1068;
    reg node1069_r;
    reg node1069_l;
    reg node1070;
    reg node1071;
    reg node1072_r;
    reg node1072_l;
    reg node1073_r;
    reg node1073_l;
    reg node1074_r;
    reg node1074_l;
    reg node1075_r;
    reg node1075_l;
    reg node1076;
    reg node1077;
    reg node1078_r;
    reg node1078_l;
    reg node1079;
    reg node1080;
    reg node1081_r;
    reg node1081_l;
    reg node1082_r;
    reg node1082_l;
    reg node1083;
    reg node1084;
    reg node1085_r;
    reg node1085_l;
    reg node1086;
    reg node1087;
    reg node1088_r;
    reg node1088_l;
    reg node1089_r;
    reg node1089_l;
    reg node1090_r;
    reg node1090_l;
    reg node1091;
    reg node1092;
    reg node1093_r;
    reg node1093_l;
    reg node1094;
    reg node1095;
    reg node1096_r;
    reg node1096_l;
    reg node1097_r;
    reg node1097_l;
    reg node1098;
    reg node1099;
    reg node1100_r;
    reg node1100_l;
    reg node1101;
    reg node1102;
    reg node1103_r;
    reg node1103_l;
    reg node1104_r;
    reg node1104_l;
    reg node1105;
    reg node1106;
    reg node1107_r;
    reg node1107_l;
    reg node1108_r;
    reg node1108_l;
    reg node1109_r;
    reg node1109_l;
    reg node1110;
    reg node1111_r;
    reg node1111_l;
    reg node1112;
    reg node1113;
    reg node1114_r;
    reg node1114_l;
    reg node1115_r;
    reg node1115_l;
    reg node1116_r;
    reg node1116_l;
    reg node1117;
    reg node1118;
    reg node1119;
    reg node1120;
    reg node1121;
    reg node1122_r;
    reg node1122_l;
    reg node1123_r;
    reg node1123_l;
    reg node1124_r;
    reg node1124_l;
    reg node1125_r;
    reg node1125_l;
    reg node1126_r;
    reg node1126_l;
    reg node1127_r;
    reg node1127_l;
    reg node1128_r;
    reg node1128_l;
    reg node1129_r;
    reg node1129_l;
    reg node1130;
    reg node1131;
    reg node1132_r;
    reg node1132_l;
    reg node1133;
    reg node1134;
    reg node1135_r;
    reg node1135_l;
    reg node1136_r;
    reg node1136_l;
    reg node1137;
    reg node1138;
    reg node1139_r;
    reg node1139_l;
    reg node1140;
    reg node1141;
    reg node1142_r;
    reg node1142_l;
    reg node1143_r;
    reg node1143_l;
    reg node1144_r;
    reg node1144_l;
    reg node1145;
    reg node1146;
    reg node1147_r;
    reg node1147_l;
    reg node1148;
    reg node1149;
    reg node1150_r;
    reg node1150_l;
    reg node1151_r;
    reg node1151_l;
    reg node1152;
    reg node1153;
    reg node1154;
    reg node1155_r;
    reg node1155_l;
    reg node1156_r;
    reg node1156_l;
    reg node1157_r;
    reg node1157_l;
    reg node1158_r;
    reg node1158_l;
    reg node1159;
    reg node1160;
    reg node1161_r;
    reg node1161_l;
    reg node1162;
    reg node1163;
    reg node1164;
    reg node1165_r;
    reg node1165_l;
    reg node1166_r;
    reg node1166_l;
    reg node1167_r;
    reg node1167_l;
    reg node1168;
    reg node1169;
    reg node1170;
    reg node1171_r;
    reg node1171_l;
    reg node1172_r;
    reg node1172_l;
    reg node1173;
    reg node1174;
    reg node1175_r;
    reg node1175_l;
    reg node1176;
    reg node1177;
    reg node1178_r;
    reg node1178_l;
    reg node1179_r;
    reg node1179_l;
    reg node1180_r;
    reg node1180_l;
    reg node1181_r;
    reg node1181_l;
    reg node1182_r;
    reg node1182_l;
    reg node1183;
    reg node1184;
    reg node1185_r;
    reg node1185_l;
    reg node1186;
    reg node1187;
    reg node1188_r;
    reg node1188_l;
    reg node1189_r;
    reg node1189_l;
    reg node1190;
    reg node1191;
    reg node1192_r;
    reg node1192_l;
    reg node1193;
    reg node1194;
    reg node1195_r;
    reg node1195_l;
    reg node1196_r;
    reg node1196_l;
    reg node1197_r;
    reg node1197_l;
    reg node1198;
    reg node1199;
    reg node1200_r;
    reg node1200_l;
    reg node1201;
    reg node1202;
    reg node1203_r;
    reg node1203_l;
    reg node1204_r;
    reg node1204_l;
    reg node1205;
    reg node1206;
    reg node1207_r;
    reg node1207_l;
    reg node1208;
    reg node1209;
    reg node1210_r;
    reg node1210_l;
    reg node1211_r;
    reg node1211_l;
    reg node1212_r;
    reg node1212_l;
    reg node1213_r;
    reg node1213_l;
    reg node1214;
    reg node1215;
    reg node1216;
    reg node1217_r;
    reg node1217_l;
    reg node1218_r;
    reg node1218_l;
    reg node1219;
    reg node1220;
    reg node1221_r;
    reg node1221_l;
    reg node1222;
    reg node1223;
    reg node1224_r;
    reg node1224_l;
    reg node1225_r;
    reg node1225_l;
    reg node1226_r;
    reg node1226_l;
    reg node1227;
    reg node1228;
    reg node1229_r;
    reg node1229_l;
    reg node1230;
    reg node1231;
    reg node1232_r;
    reg node1232_l;
    reg node1233_r;
    reg node1233_l;
    reg node1234;
    reg node1235;
    reg node1236_r;
    reg node1236_l;
    reg node1237;
    reg node1238;
    reg node1239_r;
    reg node1239_l;
    reg node1240_r;
    reg node1240_l;
    reg node1241_r;
    reg node1241_l;
    reg node1242_r;
    reg node1242_l;
    reg node1243_r;
    reg node1243_l;
    reg node1244_r;
    reg node1244_l;
    reg node1245;
    reg node1246;
    reg node1247_r;
    reg node1247_l;
    reg node1248;
    reg node1249;
    reg node1250_r;
    reg node1250_l;
    reg node1251_r;
    reg node1251_l;
    reg node1252;
    reg node1253;
    reg node1254_r;
    reg node1254_l;
    reg node1255;
    reg node1256;
    reg node1257_r;
    reg node1257_l;
    reg node1258_r;
    reg node1258_l;
    reg node1259;
    reg node1260_r;
    reg node1260_l;
    reg node1261;
    reg node1262;
    reg node1263_r;
    reg node1263_l;
    reg node1264_r;
    reg node1264_l;
    reg node1265;
    reg node1266;
    reg node1267_r;
    reg node1267_l;
    reg node1268;
    reg node1269;
    reg node1270_r;
    reg node1270_l;
    reg node1271_r;
    reg node1271_l;
    reg node1272_r;
    reg node1272_l;
    reg node1273_r;
    reg node1273_l;
    reg node1274;
    reg node1275;
    reg node1276_r;
    reg node1276_l;
    reg node1277;
    reg node1278;
    reg node1279;
    reg node1280_r;
    reg node1280_l;
    reg node1281_r;
    reg node1281_l;
    reg node1282_r;
    reg node1282_l;
    reg node1283;
    reg node1284;
    reg node1285_r;
    reg node1285_l;
    reg node1286;
    reg node1287;
    reg node1288_r;
    reg node1288_l;
    reg node1289_r;
    reg node1289_l;
    reg node1290;
    reg node1291;
    reg node1292;
    reg node1293_r;
    reg node1293_l;
    reg node1294_r;
    reg node1294_l;
    reg node1295_r;
    reg node1295_l;
    reg node1296_r;
    reg node1296_l;
    reg node1297_r;
    reg node1297_l;
    reg node1298;
    reg node1299;
    reg node1300_r;
    reg node1300_l;
    reg node1301;
    reg node1302;
    reg node1303_r;
    reg node1303_l;
    reg node1304_r;
    reg node1304_l;
    reg node1305;
    reg node1306;
    reg node1307_r;
    reg node1307_l;
    reg node1308;
    reg node1309;
    reg node1310_r;
    reg node1310_l;
    reg node1311_r;
    reg node1311_l;
    reg node1312_r;
    reg node1312_l;
    reg node1313;
    reg node1314;
    reg node1315;
    reg node1316_r;
    reg node1316_l;
    reg node1317_r;
    reg node1317_l;
    reg node1318;
    reg node1319;
    reg node1320_r;
    reg node1320_l;
    reg node1321;
    reg node1322;
    reg node1323_r;
    reg node1323_l;
    reg node1324_r;
    reg node1324_l;
    reg node1325_r;
    reg node1325_l;
    reg node1326_r;
    reg node1326_l;
    reg node1327;
    reg node1328;
    reg node1329_r;
    reg node1329_l;
    reg node1330;
    reg node1331;
    reg node1332_r;
    reg node1332_l;
    reg node1333_r;
    reg node1333_l;
    reg node1334;
    reg node1335;
    reg node1336_r;
    reg node1336_l;
    reg node1337;
    reg node1338;
    reg node1339_r;
    reg node1339_l;
    reg node1340_r;
    reg node1340_l;
    reg node1341_r;
    reg node1341_l;
    reg node1342;
    reg node1343;
    reg node1344_r;
    reg node1344_l;
    reg node1345;
    reg node1346;
    reg node1347_r;
    reg node1347_l;
    reg node1348_r;
    reg node1348_l;
    reg node1349;
    reg node1350;
    reg node1351;
    reg node1352_r;
    reg node1352_l;
    reg node1353_r;
    reg node1353_l;
    reg node1354_r;
    reg node1354_l;
    reg node1355_r;
    reg node1355_l;
    reg node1356_r;
    reg node1356_l;
    reg node1357_r;
    reg node1357_l;
    reg node1358_r;
    reg node1358_l;
    reg node1359;
    reg node1360;
    reg node1361_r;
    reg node1361_l;
    reg node1362;
    reg node1363;
    reg node1364_r;
    reg node1364_l;
    reg node1365_r;
    reg node1365_l;
    reg node1366;
    reg node1367;
    reg node1368;
    reg node1369_r;
    reg node1369_l;
    reg node1370_r;
    reg node1370_l;
    reg node1371_r;
    reg node1371_l;
    reg node1372;
    reg node1373;
    reg node1374_r;
    reg node1374_l;
    reg node1375;
    reg node1376;
    reg node1377_r;
    reg node1377_l;
    reg node1378_r;
    reg node1378_l;
    reg node1379;
    reg node1380;
    reg node1381_r;
    reg node1381_l;
    reg node1382;
    reg node1383;
    reg node1384_r;
    reg node1384_l;
    reg node1385_r;
    reg node1385_l;
    reg node1386_r;
    reg node1386_l;
    reg node1387_r;
    reg node1387_l;
    reg node1388;
    reg node1389;
    reg node1390_r;
    reg node1390_l;
    reg node1391;
    reg node1392;
    reg node1393_r;
    reg node1393_l;
    reg node1394_r;
    reg node1394_l;
    reg node1395;
    reg node1396;
    reg node1397_r;
    reg node1397_l;
    reg node1398;
    reg node1399;
    reg node1400_r;
    reg node1400_l;
    reg node1401_r;
    reg node1401_l;
    reg node1402_r;
    reg node1402_l;
    reg node1403;
    reg node1404;
    reg node1405_r;
    reg node1405_l;
    reg node1406;
    reg node1407;
    reg node1408_r;
    reg node1408_l;
    reg node1409_r;
    reg node1409_l;
    reg node1410;
    reg node1411;
    reg node1412_r;
    reg node1412_l;
    reg node1413;
    reg node1414;
    reg node1415_r;
    reg node1415_l;
    reg node1416_r;
    reg node1416_l;
    reg node1417_r;
    reg node1417_l;
    reg node1418_r;
    reg node1418_l;
    reg node1419_r;
    reg node1419_l;
    reg node1420;
    reg node1421;
    reg node1422_r;
    reg node1422_l;
    reg node1423;
    reg node1424;
    reg node1425_r;
    reg node1425_l;
    reg node1426_r;
    reg node1426_l;
    reg node1427;
    reg node1428;
    reg node1429_r;
    reg node1429_l;
    reg node1430;
    reg node1431;
    reg node1432_r;
    reg node1432_l;
    reg node1433_r;
    reg node1433_l;
    reg node1434_r;
    reg node1434_l;
    reg node1435;
    reg node1436;
    reg node1437_r;
    reg node1437_l;
    reg node1438;
    reg node1439;
    reg node1440_r;
    reg node1440_l;
    reg node1441_r;
    reg node1441_l;
    reg node1442;
    reg node1443;
    reg node1444_r;
    reg node1444_l;
    reg node1445;
    reg node1446;
    reg node1447_r;
    reg node1447_l;
    reg node1448_r;
    reg node1448_l;
    reg node1449_r;
    reg node1449_l;
    reg node1450_r;
    reg node1450_l;
    reg node1451;
    reg node1452;
    reg node1453_r;
    reg node1453_l;
    reg node1454;
    reg node1455;
    reg node1456_r;
    reg node1456_l;
    reg node1457;
    reg node1458_r;
    reg node1458_l;
    reg node1459;
    reg node1460;
    reg node1461_r;
    reg node1461_l;
    reg node1462_r;
    reg node1462_l;
    reg node1463;
    reg node1464_r;
    reg node1464_l;
    reg node1465;
    reg node1466;
    reg node1467_r;
    reg node1467_l;
    reg node1468_r;
    reg node1468_l;
    reg node1469;
    reg node1470;
    reg node1471_r;
    reg node1471_l;
    reg node1472;
    reg node1473;
    reg node1474_r;
    reg node1474_l;
    reg node1475_r;
    reg node1475_l;
    reg node1476_r;
    reg node1476_l;
    reg node1477_r;
    reg node1477_l;
    reg node1478_r;
    reg node1478_l;
    reg node1479_r;
    reg node1479_l;
    reg node1480;
    reg node1481;
    reg node1482_r;
    reg node1482_l;
    reg node1483;
    reg node1484;
    reg node1485_r;
    reg node1485_l;
    reg node1486_r;
    reg node1486_l;
    reg node1487;
    reg node1488;
    reg node1489_r;
    reg node1489_l;
    reg node1490;
    reg node1491;
    reg node1492_r;
    reg node1492_l;
    reg node1493_r;
    reg node1493_l;
    reg node1494_r;
    reg node1494_l;
    reg node1495;
    reg node1496;
    reg node1497_r;
    reg node1497_l;
    reg node1498;
    reg node1499;
    reg node1500_r;
    reg node1500_l;
    reg node1501_r;
    reg node1501_l;
    reg node1502;
    reg node1503;
    reg node1504_r;
    reg node1504_l;
    reg node1505;
    reg node1506;
    reg node1507_r;
    reg node1507_l;
    reg node1508_r;
    reg node1508_l;
    reg node1509_r;
    reg node1509_l;
    reg node1510_r;
    reg node1510_l;
    reg node1511;
    reg node1512;
    reg node1513_r;
    reg node1513_l;
    reg node1514;
    reg node1515;
    reg node1516_r;
    reg node1516_l;
    reg node1517_r;
    reg node1517_l;
    reg node1518;
    reg node1519;
    reg node1520_r;
    reg node1520_l;
    reg node1521;
    reg node1522;
    reg node1523_r;
    reg node1523_l;
    reg node1524_r;
    reg node1524_l;
    reg node1525_r;
    reg node1525_l;
    reg node1526;
    reg node1527;
    reg node1528_r;
    reg node1528_l;
    reg node1529;
    reg node1530;
    reg node1531_r;
    reg node1531_l;
    reg node1532;
    reg node1533;
    reg node1534_r;
    reg node1534_l;
    reg node1535_r;
    reg node1535_l;
    reg node1536_r;
    reg node1536_l;
    reg node1537_r;
    reg node1537_l;
    reg node1538_r;
    reg node1538_l;
    reg node1539;
    reg node1540;
    reg node1541_r;
    reg node1541_l;
    reg node1542;
    reg node1543;
    reg node1544_r;
    reg node1544_l;
    reg node1545_r;
    reg node1545_l;
    reg node1546;
    reg node1547;
    reg node1548_r;
    reg node1548_l;
    reg node1549;
    reg node1550;
    reg node1551_r;
    reg node1551_l;
    reg node1552_r;
    reg node1552_l;
    reg node1553_r;
    reg node1553_l;
    reg node1554;
    reg node1555;
    reg node1556;
    reg node1557_r;
    reg node1557_l;
    reg node1558;
    reg node1559_r;
    reg node1559_l;
    reg node1560;
    reg node1561;
    reg node1562_r;
    reg node1562_l;
    reg node1563_r;
    reg node1563_l;
    reg node1564_r;
    reg node1564_l;
    reg node1565_r;
    reg node1565_l;
    reg node1566;
    reg node1567;
    reg node1568_r;
    reg node1568_l;
    reg node1569;
    reg node1570;
    reg node1571_r;
    reg node1571_l;
    reg node1572_r;
    reg node1572_l;
    reg node1573;
    reg node1574;
    reg node1575_r;
    reg node1575_l;
    reg node1576;
    reg node1577;
    reg node1578_r;
    reg node1578_l;
    reg node1579_r;
    reg node1579_l;
    reg node1580_r;
    reg node1580_l;
    reg node1581;
    reg node1582;
    reg node1583_r;
    reg node1583_l;
    reg node1584;
    reg node1585;
    reg node1586_r;
    reg node1586_l;
    reg node1587_r;
    reg node1587_l;
    reg node1588;
    reg node1589;
    reg node1590_r;
    reg node1590_l;
    reg node1591;
    reg node1592;
    reg result0;
    reg result1;
    reg result2;
    reg result3;
    reg result4;
    reg result5;
    reg result6;
    reg result7;
    reg result8;
    reg result9;

    begin
      node0_r = pixel[429];
      node0_l = ~pixel[429];
      node1_r = node0_l & pixel[438];
      node1_l = node0_l & ~pixel[438];
      node2_r = node1_l & pixel[322];
      node2_l = node1_l & ~pixel[322];
      node3_r = node2_l & pixel[348];
      node3_l = node2_l & ~pixel[348];
      node4_r = node3_l & pixel[399];
      node4_l = node3_l & ~pixel[399];
      node5_r = node4_l & pixel[374];
      node5_l = node4_l & ~pixel[374];
      node6_r = node5_l & pixel[579];
      node6_l = node5_l & ~pixel[579];
      node7_r = node6_l & pixel[624];
      node7_l = node6_l & ~pixel[624];
      node8_r = node7_l & pixel[236];
      node8_l = node7_l & ~pixel[236];
      node9_r = node8_l & pixel[326];
      node9_l = node8_l & ~pixel[326];
      node10 = node9_l;
      node11 = node9_r;
      node12_r = node8_r & pixel[633];
      node12_l = node8_r & ~pixel[633];
      node13 = node12_l;
      node14 = node12_r;
      node15_r = node7_r & pixel[157];
      node15_l = node7_r & ~pixel[157];
      node16_r = node15_l & pixel[706];
      node16_l = node15_l & ~pixel[706];
      node17 = node16_l;
      node18 = node16_r;
      node19_r = node15_r & pixel[520];
      node19_l = node15_r & ~pixel[520];
      node20 = node19_l;
      node21 = node19_r;
      node22_r = node6_r & pixel[369];
      node22_l = node6_r & ~pixel[369];
      node23_r = node22_l & pixel[572];
      node23_l = node22_l & ~pixel[572];
      node24_r = node23_l & pixel[683];
      node24_l = node23_l & ~pixel[683];
      node25 = node24_l;
      node26 = node24_r;
      node27_r = node23_r & pixel[227];
      node27_l = node23_r & ~pixel[227];
      node28 = node27_l;
      node29 = node27_r;
      node30_r = node22_r & pixel[379];
      node30_l = node22_r & ~pixel[379];
      node31_r = node30_l & pixel[489];
      node31_l = node30_l & ~pixel[489];
      node32 = node31_l;
      node33 = node31_r;
      node34_r = node30_r & pixel[411];
      node34_l = node30_r & ~pixel[411];
      node35 = node34_l;
      node36 = node34_r;
      node37_r = node5_r & pixel[187];
      node37_l = node5_r & ~pixel[187];
      node38_r = node37_l & pixel[436];
      node38_l = node37_l & ~pixel[436];
      node39_r = node38_l & pixel[380];
      node39_l = node38_l & ~pixel[380];
      node40_r = node39_l & pixel[515];
      node40_l = node39_l & ~pixel[515];
      node41 = node40_l;
      node42 = node40_r;
      node43_r = node39_r & pixel[582];
      node43_l = node39_r & ~pixel[582];
      node44 = node43_l;
      node45 = node43_r;
      node46_r = node38_r & pixel[404];
      node46_l = node38_r & ~pixel[404];
      node47_r = node46_l & pixel[432];
      node47_l = node46_l & ~pixel[432];
      node48 = node47_l;
      node49 = node47_r;
      node50_r = node46_r & pixel[265];
      node50_l = node46_r & ~pixel[265];
      node51 = node50_l;
      node52 = node50_r;
      node53_r = node37_r & pixel[657];
      node53_l = node37_r & ~pixel[657];
      node54_r = node53_l & pixel[265];
      node54_l = node53_l & ~pixel[265];
      node55_r = node54_l & pixel[296];
      node55_l = node54_l & ~pixel[296];
      node56 = node55_l;
      node57 = node55_r;
      node58_r = node54_r & pixel[379];
      node58_l = node54_r & ~pixel[379];
      node59 = node58_l;
      node60 = node58_r;
      node61_r = node53_r & pixel[461];
      node61_l = node53_r & ~pixel[461];
      node62_r = node61_l & pixel[490];
      node62_l = node61_l & ~pixel[490];
      node63 = node62_l;
      node64 = node62_r;
      node65_r = node61_r & pixel[354];
      node65_l = node61_r & ~pixel[354];
      node66 = node65_l;
      node67 = node65_r;
      node68_r = node4_r & pixel[185];
      node68_l = node4_r & ~pixel[185];
      node69_r = node68_l & pixel[124];
      node69_l = node68_l & ~pixel[124];
      node70_r = node69_l & pixel[237];
      node70_l = node69_l & ~pixel[237];
      node71_r = node70_l & pixel[188];
      node71_l = node70_l & ~pixel[188];
      node72_r = node71_l & pixel[575];
      node72_l = node71_l & ~pixel[575];
      node73 = node72_l;
      node74 = node72_r;
      node75_r = node71_r & pixel[408];
      node75_l = node71_r & ~pixel[408];
      node76 = node75_l;
      node77 = node75_r;
      node78_r = node70_r & pixel[568];
      node78_l = node70_r & ~pixel[568];
      node79_r = node78_l & pixel[414];
      node79_l = node78_l & ~pixel[414];
      node80 = node79_l;
      node81 = node79_r;
      node82_r = node78_r & pixel[490];
      node82_l = node78_r & ~pixel[490];
      node83 = node82_l;
      node84 = node82_r;
      node85_r = node69_r & pixel[408];
      node85_l = node69_r & ~pixel[408];
      node86_r = node85_l & pixel[629];
      node86_l = node85_l & ~pixel[629];
      node87_r = node86_l & pixel[207];
      node87_l = node86_l & ~pixel[207];
      node88 = node87_l;
      node89 = node87_r;
      node90_r = node86_r & pixel[435];
      node90_l = node86_r & ~pixel[435];
      node91 = node90_l;
      node92 = node90_r;
      node93_r = node85_r & pixel[315];
      node93_l = node85_r & ~pixel[315];
      node94_r = node93_l & pixel[324];
      node94_l = node93_l & ~pixel[324];
      node95 = node94_l;
      node96 = node94_r;
      node97 = node93_r;
      node98_r = node68_r & pixel[408];
      node98_l = node68_r & ~pixel[408];
      node99_r = node98_l & pixel[714];
      node99_l = node98_l & ~pixel[714];
      node100_r = node99_l & pixel[221];
      node100_l = node99_l & ~pixel[221];
      node101_r = node100_l & pixel[261];
      node101_l = node100_l & ~pixel[261];
      node102 = node101_l;
      node103 = node101_r;
      node104 = node100_r;
      node105 = node99_r;
      node106_r = node98_r & pixel[101];
      node106_l = node98_r & ~pixel[101];
      node107_r = node106_l & pixel[273];
      node107_l = node106_l & ~pixel[273];
      node108_r = node107_l & pixel[499];
      node108_l = node107_l & ~pixel[499];
      node109 = node108_l;
      node110 = node108_r;
      node111_r = node107_r & pixel[597];
      node111_l = node107_r & ~pixel[597];
      node112 = node111_l;
      node113 = node111_r;
      node114 = node106_r;
      node115_r = node3_r & pixel[407];
      node115_l = node3_r & ~pixel[407];
      node116_r = node115_l & pixel[360];
      node116_l = node115_l & ~pixel[360];
      node117_r = node116_l & pixel[626];
      node117_l = node116_l & ~pixel[626];
      node118_r = node117_l & pixel[550];
      node118_l = node117_l & ~pixel[550];
      node119_r = node118_l & pixel[381];
      node119_l = node118_l & ~pixel[381];
      node120_r = node119_l & pixel[657];
      node120_l = node119_l & ~pixel[657];
      node121 = node120_l;
      node122 = node120_r;
      node123_r = node119_r & pixel[572];
      node123_l = node119_r & ~pixel[572];
      node124 = node123_l;
      node125 = node123_r;
      node126_r = node118_r & pixel[544];
      node126_l = node118_r & ~pixel[544];
      node127_r = node126_l & pixel[263];
      node127_l = node126_l & ~pixel[263];
      node128 = node127_l;
      node129 = node127_r;
      node130_r = node126_r & pixel[543];
      node130_l = node126_r & ~pixel[543];
      node131 = node130_l;
      node132 = node130_r;
      node133_r = node117_r & pixel[426];
      node133_l = node117_r & ~pixel[426];
      node134_r = node133_l & pixel[375];
      node134_l = node133_l & ~pixel[375];
      node135_r = node134_l & pixel[295];
      node135_l = node134_l & ~pixel[295];
      node136 = node135_l;
      node137 = node135_r;
      node138_r = node134_r & pixel[218];
      node138_l = node134_r & ~pixel[218];
      node139 = node138_l;
      node140 = node138_r;
      node141_r = node133_r & pixel[274];
      node141_l = node133_r & ~pixel[274];
      node142_r = node141_l & pixel[403];
      node142_l = node141_l & ~pixel[403];
      node143 = node142_l;
      node144 = node142_r;
      node145_r = node141_r & pixel[358];
      node145_l = node141_r & ~pixel[358];
      node146 = node145_l;
      node147 = node145_r;
      node148 = node116_r;
      node149_r = node115_r & pixel[488];
      node149_l = node115_r & ~pixel[488];
      node150_r = node149_l & pixel[326];
      node150_l = node149_l & ~pixel[326];
      node151_r = node150_l & pixel[627];
      node151_l = node150_l & ~pixel[627];
      node152_r = node151_l & pixel[541];
      node152_l = node151_l & ~pixel[541];
      node153_r = node152_l & pixel[352];
      node153_l = node152_l & ~pixel[352];
      node154 = node153_l;
      node155 = node153_r;
      node156_r = node152_r & pixel[299];
      node156_l = node152_r & ~pixel[299];
      node157 = node156_l;
      node158 = node156_r;
      node159_r = node151_r & pixel[425];
      node159_l = node151_r & ~pixel[425];
      node160_r = node159_l & pixel[134];
      node160_l = node159_l & ~pixel[134];
      node161 = node160_l;
      node162 = node160_r;
      node163_r = node159_r & pixel[343];
      node163_l = node159_r & ~pixel[343];
      node164 = node163_l;
      node165 = node163_r;
      node166_r = node150_r & pixel[660];
      node166_l = node150_r & ~pixel[660];
      node167_r = node166_l & pixel[153];
      node167_l = node166_l & ~pixel[153];
      node168_r = node167_l & pixel[565];
      node168_l = node167_l & ~pixel[565];
      node169 = node168_l;
      node170 = node168_r;
      node171_r = node167_r & pixel[373];
      node171_l = node167_r & ~pixel[373];
      node172 = node171_l;
      node173 = node171_r;
      node174_r = node166_r & pixel[319];
      node174_l = node166_r & ~pixel[319];
      node175_r = node174_l & pixel[466];
      node175_l = node174_l & ~pixel[466];
      node176 = node175_l;
      node177 = node175_r;
      node178_r = node174_r & pixel[656];
      node178_l = node174_r & ~pixel[656];
      node179 = node178_l;
      node180 = node178_r;
      node181_r = node149_r & pixel[405];
      node181_l = node149_r & ~pixel[405];
      node182_r = node181_l & pixel[598];
      node182_l = node181_l & ~pixel[598];
      node183_r = node182_l & pixel[656];
      node183_l = node182_l & ~pixel[656];
      node184_r = node183_l & pixel[686];
      node184_l = node183_l & ~pixel[686];
      node185 = node184_l;
      node186 = node184_r;
      node187_r = node183_r & pixel[624];
      node187_l = node183_r & ~pixel[624];
      node188 = node187_l;
      node189 = node187_r;
      node190_r = node182_r & pixel[709];
      node190_l = node182_r & ~pixel[709];
      node191_r = node190_l & pixel[707];
      node191_l = node190_l & ~pixel[707];
      node192 = node191_l;
      node193 = node191_r;
      node194 = node190_r;
      node195_r = node181_r & pixel[186];
      node195_l = node181_r & ~pixel[186];
      node196_r = node195_l & pixel[270];
      node196_l = node195_l & ~pixel[270];
      node197_r = node196_l & pixel[184];
      node197_l = node196_l & ~pixel[184];
      node198 = node197_l;
      node199 = node197_r;
      node200_r = node196_r & pixel[632];
      node200_l = node196_r & ~pixel[632];
      node201 = node200_l;
      node202 = node200_r;
      node203_r = node195_r & pixel[656];
      node203_l = node195_r & ~pixel[656];
      node204_r = node203_l & pixel[487];
      node204_l = node203_l & ~pixel[487];
      node205 = node204_l;
      node206 = node204_r;
      node207_r = node203_r & pixel[626];
      node207_l = node203_r & ~pixel[626];
      node208 = node207_l;
      node209 = node207_r;
      node210_r = node2_r & pixel[550];
      node210_l = node2_r & ~pixel[550];
      node211_r = node210_l & pixel[347];
      node211_l = node210_l & ~pixel[347];
      node212_r = node211_l & pixel[218];
      node212_l = node211_l & ~pixel[218];
      node213_r = node212_l & pixel[272];
      node213_l = node212_l & ~pixel[272];
      node214_r = node213_l & pixel[517];
      node214_l = node213_l & ~pixel[517];
      node215_r = node214_l & pixel[157];
      node215_l = node214_l & ~pixel[157];
      node216_r = node215_l & pixel[656];
      node216_l = node215_l & ~pixel[656];
      node217 = node216_l;
      node218 = node216_r;
      node219_r = node215_r & pixel[460];
      node219_l = node215_r & ~pixel[460];
      node220 = node219_l;
      node221 = node219_r;
      node222_r = node214_r & pixel[176];
      node222_l = node214_r & ~pixel[176];
      node223_r = node222_l & pixel[291];
      node223_l = node222_l & ~pixel[291];
      node224 = node223_l;
      node225 = node223_r;
      node226_r = node222_r & pixel[634];
      node226_l = node222_r & ~pixel[634];
      node227 = node226_l;
      node228 = node226_r;
      node229_r = node213_r & pixel[657];
      node229_l = node213_r & ~pixel[657];
      node230_r = node229_l & pixel[602];
      node230_l = node229_l & ~pixel[602];
      node231_r = node230_l & pixel[624];
      node231_l = node230_l & ~pixel[624];
      node232 = node231_l;
      node233 = node231_r;
      node234_r = node230_r & pixel[471];
      node234_l = node230_r & ~pixel[471];
      node235 = node234_l;
      node236 = node234_r;
      node237_r = node229_r & pixel[738];
      node237_l = node229_r & ~pixel[738];
      node238_r = node237_l & pixel[343];
      node238_l = node237_l & ~pixel[343];
      node239 = node238_l;
      node240 = node238_r;
      node241 = node237_r;
      node242_r = node212_r & pixel[600];
      node242_l = node212_r & ~pixel[600];
      node243_r = node242_l & pixel[683];
      node243_l = node242_l & ~pixel[683];
      node244_r = node243_l & pixel[519];
      node244_l = node243_l & ~pixel[519];
      node245_r = node244_l & pixel[541];
      node245_l = node244_l & ~pixel[541];
      node246 = node245_l;
      node247 = node245_r;
      node248_r = node244_r & pixel[517];
      node248_l = node244_r & ~pixel[517];
      node249 = node248_l;
      node250 = node248_r;
      node251_r = node243_r & pixel[415];
      node251_l = node243_r & ~pixel[415];
      node252_r = node251_l & pixel[157];
      node252_l = node251_l & ~pixel[157];
      node253 = node252_l;
      node254 = node252_r;
      node255 = node251_r;
      node256_r = node242_r & pixel[273];
      node256_l = node242_r & ~pixel[273];
      node257_r = node256_l & pixel[520];
      node257_l = node256_l & ~pixel[520];
      node258_r = node257_l & pixel[488];
      node258_l = node257_l & ~pixel[488];
      node259 = node258_l;
      node260 = node258_r;
      node261_r = node257_r & pixel[355];
      node261_l = node257_r & ~pixel[355];
      node262 = node261_l;
      node263 = node261_r;
      node264_r = node256_r & pixel[354];
      node264_l = node256_r & ~pixel[354];
      node265_r = node264_l & pixel[331];
      node265_l = node264_l & ~pixel[331];
      node266 = node265_l;
      node267 = node265_r;
      node268_r = node264_r & pixel[182];
      node268_l = node264_r & ~pixel[182];
      node269 = node268_l;
      node270 = node268_r;
      node271_r = node211_r & pixel[510];
      node271_l = node211_r & ~pixel[510];
      node272_r = node271_l & pixel[597];
      node272_l = node271_l & ~pixel[597];
      node273_r = node272_l & pixel[153];
      node273_l = node272_l & ~pixel[153];
      node274_r = node273_l & pixel[379];
      node274_l = node273_l & ~pixel[379];
      node275_r = node274_l & pixel[409];
      node275_l = node274_l & ~pixel[409];
      node276 = node275_l;
      node277 = node275_r;
      node278_r = node274_r & pixel[211];
      node278_l = node274_r & ~pixel[211];
      node279 = node278_l;
      node280 = node278_r;
      node281_r = node273_r & pixel[518];
      node281_l = node273_r & ~pixel[518];
      node282_r = node281_l & pixel[319];
      node282_l = node281_l & ~pixel[319];
      node283 = node282_l;
      node284 = node282_r;
      node285_r = node281_r & pixel[292];
      node285_l = node281_r & ~pixel[292];
      node286 = node285_l;
      node287 = node285_r;
      node288_r = node272_r & pixel[353];
      node288_l = node272_r & ~pixel[353];
      node289_r = node288_l & pixel[596];
      node289_l = node288_l & ~pixel[596];
      node290_r = node289_l & pixel[208];
      node290_l = node289_l & ~pixel[208];
      node291 = node290_l;
      node292 = node290_r;
      node293_r = node289_r & pixel[203];
      node293_l = node289_r & ~pixel[203];
      node294 = node293_l;
      node295 = node293_r;
      node296_r = node288_r & pixel[441];
      node296_l = node288_r & ~pixel[441];
      node297_r = node296_l & pixel[514];
      node297_l = node296_l & ~pixel[514];
      node298 = node297_l;
      node299 = node297_r;
      node300_r = node296_r & pixel[261];
      node300_l = node296_r & ~pixel[261];
      node301 = node300_l;
      node302 = node300_r;
      node303_r = node271_r & pixel[579];
      node303_l = node271_r & ~pixel[579];
      node304_r = node303_l & pixel[126];
      node304_l = node303_l & ~pixel[126];
      node305_r = node304_l & pixel[650];
      node305_l = node304_l & ~pixel[650];
      node306_r = node305_l & pixel[293];
      node306_l = node305_l & ~pixel[293];
      node307 = node306_l;
      node308 = node306_r;
      node309_r = node305_r & pixel[354];
      node309_l = node305_r & ~pixel[354];
      node310 = node309_l;
      node311 = node309_r;
      node312_r = node304_r & pixel[383];
      node312_l = node304_r & ~pixel[383];
      node313 = node312_l;
      node314 = node312_r;
      node315_r = node303_r & pixel[158];
      node315_l = node303_r & ~pixel[158];
      node316_r = node315_l & pixel[148];
      node316_l = node315_l & ~pixel[148];
      node317_r = node316_l & pixel[381];
      node317_l = node316_l & ~pixel[381];
      node318 = node317_l;
      node319 = node317_r;
      node320_r = node316_r & pixel[582];
      node320_l = node316_r & ~pixel[582];
      node321 = node320_l;
      node322 = node320_r;
      node323_r = node315_r & pixel[376];
      node323_l = node315_r & ~pixel[376];
      node324 = node323_l;
      node325_r = node323_r & pixel[177];
      node325_l = node323_r & ~pixel[177];
      node326 = node325_l;
      node327 = node325_r;
      node328_r = node210_r & pixel[555];
      node328_l = node210_r & ~pixel[555];
      node329_r = node328_l & pixel[482];
      node329_l = node328_l & ~pixel[482];
      node330_r = node329_l & pixel[459];
      node330_l = node329_l & ~pixel[459];
      node331_r = node330_l & pixel[517];
      node331_l = node330_l & ~pixel[517];
      node332_r = node331_l & pixel[404];
      node332_l = node331_l & ~pixel[404];
      node333_r = node332_l & pixel[629];
      node333_l = node332_l & ~pixel[629];
      node334 = node333_l;
      node335 = node333_r;
      node336_r = node332_r & pixel[289];
      node336_l = node332_r & ~pixel[289];
      node337 = node336_l;
      node338 = node336_r;
      node339_r = node331_r & pixel[660];
      node339_l = node331_r & ~pixel[660];
      node340_r = node339_l & pixel[266];
      node340_l = node339_l & ~pixel[266];
      node341 = node340_l;
      node342 = node340_r;
      node343_r = node339_r & pixel[347];
      node343_l = node339_r & ~pixel[347];
      node344 = node343_l;
      node345 = node343_r;
      node346_r = node330_r & pixel[262];
      node346_l = node330_r & ~pixel[262];
      node347_r = node346_l & pixel[103];
      node347_l = node346_l & ~pixel[103];
      node348_r = node347_l & pixel[552];
      node348_l = node347_l & ~pixel[552];
      node349 = node348_l;
      node350 = node348_r;
      node351_r = node347_r & pixel[626];
      node351_l = node347_r & ~pixel[626];
      node352 = node351_l;
      node353 = node351_r;
      node354_r = node346_r & pixel[318];
      node354_l = node346_r & ~pixel[318];
      node355_r = node354_l & pixel[544];
      node355_l = node354_l & ~pixel[544];
      node356 = node355_l;
      node357 = node355_r;
      node358_r = node354_r & pixel[610];
      node358_l = node354_r & ~pixel[610];
      node359 = node358_l;
      node360 = node358_r;
      node361_r = node329_r & pixel[370];
      node361_l = node329_r & ~pixel[370];
      node362_r = node361_l & pixel[330];
      node362_l = node361_l & ~pixel[330];
      node363_r = node362_l & pixel[247];
      node363_l = node362_l & ~pixel[247];
      node364_r = node363_l & pixel[458];
      node364_l = node363_l & ~pixel[458];
      node365 = node364_l;
      node366 = node364_r;
      node367_r = node363_r & pixel[128];
      node367_l = node363_r & ~pixel[128];
      node368 = node367_l;
      node369 = node367_r;
      node370_r = node362_r & pixel[292];
      node370_l = node362_r & ~pixel[292];
      node371_r = node370_l & pixel[406];
      node371_l = node370_l & ~pixel[406];
      node372 = node371_l;
      node373 = node371_r;
      node374 = node370_r;
      node375_r = node361_r & pixel[460];
      node375_l = node361_r & ~pixel[460];
      node376_r = node375_l & pixel[717];
      node376_l = node375_l & ~pixel[717];
      node377_r = node376_l & pixel[148];
      node377_l = node376_l & ~pixel[148];
      node378 = node377_l;
      node379 = node377_r;
      node380 = node376_r;
      node381 = node375_r;
      node382_r = node328_r & pixel[331];
      node382_l = node328_r & ~pixel[331];
      node383_r = node382_l & pixel[415];
      node383_l = node382_l & ~pixel[415];
      node384_r = node383_l & pixel[488];
      node384_l = node383_l & ~pixel[488];
      node385_r = node384_l & pixel[557];
      node385_l = node384_l & ~pixel[557];
      node386_r = node385_l & pixel[435];
      node386_l = node385_l & ~pixel[435];
      node387 = node386_l;
      node388 = node386_r;
      node389_r = node385_r & pixel[266];
      node389_l = node385_r & ~pixel[266];
      node390 = node389_l;
      node391 = node389_r;
      node392 = node384_r;
      node393_r = node383_r & pixel[157];
      node393_l = node383_r & ~pixel[157];
      node394_r = node393_l & pixel[456];
      node394_l = node393_l & ~pixel[456];
      node395_r = node394_l & pixel[605];
      node395_l = node394_l & ~pixel[605];
      node396 = node395_l;
      node397 = node395_r;
      node398_r = node394_r & pixel[240];
      node398_l = node394_r & ~pixel[240];
      node399 = node398_l;
      node400 = node398_r;
      node401_r = node393_r & pixel[208];
      node401_l = node393_r & ~pixel[208];
      node402 = node401_l;
      node403_r = node401_r & pixel[315];
      node403_l = node401_r & ~pixel[315];
      node404 = node403_l;
      node405 = node403_r;
      node406_r = node382_r & pixel[633];
      node406_l = node382_r & ~pixel[633];
      node407 = node406_l;
      node408 = node406_r;
      node409_r = node1_r & pixel[180];
      node409_l = node1_r & ~pixel[180];
      node410_r = node409_l & pixel[287];
      node410_l = node409_l & ~pixel[287];
      node411_r = node410_l & pixel[431];
      node411_l = node410_l & ~pixel[431];
      node412_r = node411_l & pixel[568];
      node412_l = node411_l & ~pixel[568];
      node413_r = node412_l & pixel[350];
      node413_l = node412_l & ~pixel[350];
      node414_r = node413_l & pixel[483];
      node414_l = node413_l & ~pixel[483];
      node415_r = node414_l & pixel[269];
      node415_l = node414_l & ~pixel[269];
      node416_r = node415_l & pixel[432];
      node416_l = node415_l & ~pixel[432];
      node417 = node416_l;
      node418 = node416_r;
      node419_r = node415_r & pixel[593];
      node419_l = node415_r & ~pixel[593];
      node420 = node419_l;
      node421 = node419_r;
      node422_r = node414_r & pixel[355];
      node422_l = node414_r & ~pixel[355];
      node423_r = node422_l & pixel[651];
      node423_l = node422_l & ~pixel[651];
      node424 = node423_l;
      node425 = node423_r;
      node426_r = node422_r & pixel[317];
      node426_l = node422_r & ~pixel[317];
      node427 = node426_l;
      node428 = node426_r;
      node429_r = node413_r & pixel[522];
      node429_l = node413_r & ~pixel[522];
      node430_r = node429_l & pixel[370];
      node430_l = node429_l & ~pixel[370];
      node431_r = node430_l & pixel[607];
      node431_l = node430_l & ~pixel[607];
      node432 = node431_l;
      node433 = node431_r;
      node434_r = node430_r & pixel[608];
      node434_l = node430_r & ~pixel[608];
      node435 = node434_l;
      node436 = node434_r;
      node437_r = node429_r & pixel[291];
      node437_l = node429_r & ~pixel[291];
      node438_r = node437_l & pixel[379];
      node438_l = node437_l & ~pixel[379];
      node439 = node438_l;
      node440 = node438_r;
      node441_r = node437_r & pixel[328];
      node441_l = node437_r & ~pixel[328];
      node442 = node441_l;
      node443 = node441_r;
      node444_r = node412_r & pixel[219];
      node444_l = node412_r & ~pixel[219];
      node445_r = node444_l & pixel[514];
      node445_l = node444_l & ~pixel[514];
      node446_r = node445_l & pixel[330];
      node446_l = node445_l & ~pixel[330];
      node447_r = node446_l & pixel[126];
      node447_l = node446_l & ~pixel[126];
      node448 = node447_l;
      node449 = node447_r;
      node450_r = node446_r & pixel[406];
      node450_l = node446_r & ~pixel[406];
      node451 = node450_l;
      node452 = node450_r;
      node453_r = node445_r & pixel[291];
      node453_l = node445_r & ~pixel[291];
      node454_r = node453_l & pixel[294];
      node454_l = node453_l & ~pixel[294];
      node455 = node454_l;
      node456 = node454_r;
      node457_r = node453_r & pixel[328];
      node457_l = node453_r & ~pixel[328];
      node458 = node457_l;
      node459 = node457_r;
      node460_r = node444_r & pixel[441];
      node460_l = node444_r & ~pixel[441];
      node461_r = node460_l & pixel[735];
      node461_l = node460_l & ~pixel[735];
      node462_r = node461_l & pixel[384];
      node462_l = node461_l & ~pixel[384];
      node463 = node462_l;
      node464 = node462_r;
      node465 = node461_r;
      node466_r = node460_r & pixel[522];
      node466_l = node460_r & ~pixel[522];
      node467 = node466_l;
      node468_r = node466_r & pixel[344];
      node468_l = node466_r & ~pixel[344];
      node469 = node468_l;
      node470 = node468_r;
      node471_r = node411_r & pixel[514];
      node471_l = node411_r & ~pixel[514];
      node472_r = node471_l & pixel[355];
      node472_l = node471_l & ~pixel[355];
      node473_r = node472_l & pixel[596];
      node473_l = node472_l & ~pixel[596];
      node474_r = node473_l & pixel[544];
      node474_l = node473_l & ~pixel[544];
      node475_r = node474_l & pixel[716];
      node475_l = node474_l & ~pixel[716];
      node476 = node475_l;
      node477 = node475_r;
      node478_r = node474_r & pixel[270];
      node478_l = node474_r & ~pixel[270];
      node479 = node478_l;
      node480 = node478_r;
      node481_r = node473_r & pixel[325];
      node481_l = node473_r & ~pixel[325];
      node482_r = node481_l & pixel[203];
      node482_l = node481_l & ~pixel[203];
      node483 = node482_l;
      node484 = node482_r;
      node485_r = node481_r & pixel[249];
      node485_l = node481_r & ~pixel[249];
      node486 = node485_l;
      node487 = node485_r;
      node488_r = node472_r & pixel[564];
      node488_l = node472_r & ~pixel[564];
      node489_r = node488_l & pixel[211];
      node489_l = node488_l & ~pixel[211];
      node490_r = node489_l & pixel[121];
      node490_l = node489_l & ~pixel[121];
      node491 = node490_l;
      node492 = node490_r;
      node493_r = node489_r & pixel[400];
      node493_l = node489_r & ~pixel[400];
      node494 = node493_l;
      node495 = node493_r;
      node496_r = node488_r & pixel[489];
      node496_l = node488_r & ~pixel[489];
      node497_r = node496_l & pixel[182];
      node497_l = node496_l & ~pixel[182];
      node498 = node497_l;
      node499 = node497_r;
      node500 = node496_r;
      node501_r = node471_r & pixel[297];
      node501_l = node471_r & ~pixel[297];
      node502_r = node501_l & pixel[356];
      node502_l = node501_l & ~pixel[356];
      node503_r = node502_l & pixel[301];
      node503_l = node502_l & ~pixel[301];
      node504_r = node503_l & pixel[416];
      node504_l = node503_l & ~pixel[416];
      node505 = node504_l;
      node506 = node504_r;
      node507_r = node503_r & pixel[485];
      node507_l = node503_r & ~pixel[485];
      node508 = node507_l;
      node509 = node507_r;
      node510_r = node502_r & pixel[509];
      node510_l = node502_r & ~pixel[509];
      node511_r = node510_l & pixel[303];
      node511_l = node510_l & ~pixel[303];
      node512 = node511_l;
      node513 = node511_r;
      node514_r = node510_r & pixel[566];
      node514_l = node510_r & ~pixel[566];
      node515 = node514_l;
      node516 = node514_r;
      node517_r = node501_r & pixel[264];
      node517_l = node501_r & ~pixel[264];
      node518_r = node517_l & pixel[322];
      node518_l = node517_l & ~pixel[322];
      node519_r = node518_l & pixel[288];
      node519_l = node518_l & ~pixel[288];
      node520 = node519_l;
      node521 = node519_r;
      node522_r = node518_r & pixel[458];
      node522_l = node518_r & ~pixel[458];
      node523 = node522_l;
      node524 = node522_r;
      node525_r = node517_r & pixel[623];
      node525_l = node517_r & ~pixel[623];
      node526_r = node525_l & pixel[218];
      node526_l = node525_l & ~pixel[218];
      node527 = node526_l;
      node528 = node526_r;
      node529_r = node525_r & pixel[526];
      node529_l = node525_r & ~pixel[526];
      node530 = node529_l;
      node531 = node529_r;
      node532_r = node410_r & pixel[461];
      node532_l = node410_r & ~pixel[461];
      node533_r = node532_l & pixel[401];
      node533_l = node532_l & ~pixel[401];
      node534_r = node533_l & pixel[510];
      node534_l = node533_l & ~pixel[510];
      node535_r = node534_l & pixel[403];
      node535_l = node534_l & ~pixel[403];
      node536_r = node535_l & pixel[459];
      node536_l = node535_l & ~pixel[459];
      node537_r = node536_l & pixel[405];
      node537_l = node536_l & ~pixel[405];
      node538 = node537_l;
      node539 = node537_r;
      node540_r = node536_r & pixel[661];
      node540_l = node536_r & ~pixel[661];
      node541 = node540_l;
      node542 = node540_r;
      node543_r = node535_r & pixel[464];
      node543_l = node535_r & ~pixel[464];
      node544 = node543_l;
      node545_r = node543_r & pixel[657];
      node545_l = node543_r & ~pixel[657];
      node546 = node545_l;
      node547 = node545_r;
      node548_r = node534_r & pixel[491];
      node548_l = node534_r & ~pixel[491];
      node549_r = node548_l & pixel[540];
      node549_l = node548_l & ~pixel[540];
      node550_r = node549_l & pixel[220];
      node550_l = node549_l & ~pixel[220];
      node551 = node550_l;
      node552 = node550_r;
      node553_r = node549_r & pixel[575];
      node553_l = node549_r & ~pixel[575];
      node554 = node553_l;
      node555 = node553_r;
      node556_r = node548_r & pixel[262];
      node556_l = node548_r & ~pixel[262];
      node557_r = node556_l & pixel[257];
      node557_l = node556_l & ~pixel[257];
      node558 = node557_l;
      node559 = node557_r;
      node560 = node556_r;
      node561_r = node533_r & pixel[378];
      node561_l = node533_r & ~pixel[378];
      node562_r = node561_l & pixel[513];
      node562_l = node561_l & ~pixel[513];
      node563_r = node562_l & pixel[317];
      node563_l = node562_l & ~pixel[317];
      node564_r = node563_l & pixel[213];
      node564_l = node563_l & ~pixel[213];
      node565 = node564_l;
      node566 = node564_r;
      node567_r = node563_r & pixel[230];
      node567_l = node563_r & ~pixel[230];
      node568 = node567_l;
      node569 = node567_r;
      node570_r = node562_r & pixel[633];
      node570_l = node562_r & ~pixel[633];
      node571_r = node570_l & pixel[66];
      node571_l = node570_l & ~pixel[66];
      node572 = node571_l;
      node573 = node571_r;
      node574 = node570_r;
      node575_r = node561_r & pixel[217];
      node575_l = node561_r & ~pixel[217];
      node576_r = node575_l & pixel[237];
      node576_l = node575_l & ~pixel[237];
      node577_r = node576_l & pixel[274];
      node577_l = node576_l & ~pixel[274];
      node578 = node577_l;
      node579 = node577_r;
      node580_r = node576_r & pixel[368];
      node580_l = node576_r & ~pixel[368];
      node581 = node580_l;
      node582 = node580_r;
      node583_r = node575_r & pixel[657];
      node583_l = node575_r & ~pixel[657];
      node584_r = node583_l & pixel[211];
      node584_l = node583_l & ~pixel[211];
      node585 = node584_l;
      node586 = node584_r;
      node587_r = node583_r & pixel[239];
      node587_l = node583_r & ~pixel[239];
      node588 = node587_l;
      node589 = node587_r;
      node590_r = node532_r & pixel[656];
      node590_l = node532_r & ~pixel[656];
      node591_r = node590_l & pixel[264];
      node591_l = node590_l & ~pixel[264];
      node592_r = node591_l & pixel[209];
      node592_l = node591_l & ~pixel[209];
      node593_r = node592_l & pixel[653];
      node593_l = node592_l & ~pixel[653];
      node594_r = node593_l & pixel[427];
      node594_l = node593_l & ~pixel[427];
      node595 = node594_l;
      node596 = node594_r;
      node597 = node593_r;
      node598_r = node592_r & pixel[398];
      node598_l = node592_r & ~pixel[398];
      node599_r = node598_l & pixel[208];
      node599_l = node598_l & ~pixel[208];
      node600 = node599_l;
      node601 = node599_r;
      node602 = node598_r;
      node603_r = node591_r & pixel[456];
      node603_l = node591_r & ~pixel[456];
      node604_r = node603_l & pixel[707];
      node604_l = node603_l & ~pixel[707];
      node605_r = node604_l & pixel[527];
      node605_l = node604_l & ~pixel[527];
      node606 = node605_l;
      node607 = node605_r;
      node608_r = node604_r & pixel[572];
      node608_l = node604_r & ~pixel[572];
      node609 = node608_l;
      node610 = node608_r;
      node611_r = node603_r & pixel[599];
      node611_l = node603_r & ~pixel[599];
      node612_r = node611_l & pixel[356];
      node612_l = node611_l & ~pixel[356];
      node613 = node612_l;
      node614 = node612_r;
      node615_r = node611_r & pixel[294];
      node615_l = node611_r & ~pixel[294];
      node616 = node615_l;
      node617 = node615_r;
      node618_r = node590_r & pixel[376];
      node618_l = node590_r & ~pixel[376];
      node619_r = node618_l & pixel[480];
      node619_l = node618_l & ~pixel[480];
      node620_r = node619_l & pixel[456];
      node620_l = node619_l & ~pixel[456];
      node621_r = node620_l & pixel[149];
      node621_l = node620_l & ~pixel[149];
      node622 = node621_l;
      node623 = node621_r;
      node624_r = node620_r & pixel[631];
      node624_l = node620_r & ~pixel[631];
      node625 = node624_l;
      node626 = node624_r;
      node627 = node619_r;
      node628_r = node618_r & pixel[657];
      node628_l = node618_r & ~pixel[657];
      node629_r = node628_l & pixel[190];
      node629_l = node628_l & ~pixel[190];
      node630 = node629_l;
      node631 = node629_r;
      node632_r = node628_r & pixel[540];
      node632_l = node628_r & ~pixel[540];
      node633_r = node632_l & pixel[712];
      node633_l = node632_l & ~pixel[712];
      node634 = node633_l;
      node635 = node633_r;
      node636 = node632_r;
      node637_r = node409_r & pixel[351];
      node637_l = node409_r & ~pixel[351];
      node638_r = node637_l & pixel[404];
      node638_l = node637_l & ~pixel[404];
      node639_r = node638_l & pixel[514];
      node639_l = node638_l & ~pixel[514];
      node640_r = node639_l & pixel[709];
      node640_l = node639_l & ~pixel[709];
      node641_r = node640_l & pixel[712];
      node641_l = node640_l & ~pixel[712];
      node642_r = node641_l & pixel[454];
      node642_l = node641_l & ~pixel[454];
      node643_r = node642_l & pixel[573];
      node643_l = node642_l & ~pixel[573];
      node644 = node643_l;
      node645 = node643_r;
      node646_r = node642_r & pixel[651];
      node646_l = node642_r & ~pixel[651];
      node647 = node646_l;
      node648 = node646_r;
      node649_r = node641_r & pixel[546];
      node649_l = node641_r & ~pixel[546];
      node650_r = node649_l & pixel[260];
      node650_l = node649_l & ~pixel[260];
      node651 = node650_l;
      node652 = node650_r;
      node653_r = node649_r & pixel[512];
      node653_l = node649_r & ~pixel[512];
      node654 = node653_l;
      node655 = node653_r;
      node656_r = node640_r & pixel[285];
      node656_l = node640_r & ~pixel[285];
      node657_r = node656_l & pixel[349];
      node657_l = node656_l & ~pixel[349];
      node658 = node657_l;
      node659_r = node657_r & pixel[373];
      node659_l = node657_r & ~pixel[373];
      node660 = node659_l;
      node661 = node659_r;
      node662_r = node656_r & pixel[370];
      node662_l = node656_r & ~pixel[370];
      node663_r = node662_l & pixel[258];
      node663_l = node662_l & ~pixel[258];
      node664 = node663_l;
      node665 = node663_r;
      node666 = node662_r;
      node667_r = node639_r & pixel[691];
      node667_l = node639_r & ~pixel[691];
      node668_r = node667_l & pixel[572];
      node668_l = node667_l & ~pixel[572];
      node669_r = node668_l & pixel[184];
      node669_l = node668_l & ~pixel[184];
      node670_r = node669_l & pixel[400];
      node670_l = node669_l & ~pixel[400];
      node671 = node670_l;
      node672 = node670_r;
      node673_r = node669_r & pixel[597];
      node673_l = node669_r & ~pixel[597];
      node674 = node673_l;
      node675 = node673_r;
      node676_r = node668_r & pixel[270];
      node676_l = node668_r & ~pixel[270];
      node677_r = node676_l & pixel[624];
      node677_l = node676_l & ~pixel[624];
      node678 = node677_l;
      node679 = node677_r;
      node680_r = node676_r & pixel[399];
      node680_l = node676_r & ~pixel[399];
      node681 = node680_l;
      node682 = node680_r;
      node683_r = node667_r & pixel[202];
      node683_l = node667_r & ~pixel[202];
      node684_r = node683_l & pixel[371];
      node684_l = node683_l & ~pixel[371];
      node685_r = node684_l & pixel[370];
      node685_l = node684_l & ~pixel[370];
      node686 = node685_l;
      node687 = node685_r;
      node688_r = node684_r & pixel[192];
      node688_l = node684_r & ~pixel[192];
      node689 = node688_l;
      node690 = node688_r;
      node691_r = node683_r & pixel[555];
      node691_l = node683_r & ~pixel[555];
      node692 = node691_l;
      node693 = node691_r;
      node694_r = node638_r & pixel[382];
      node694_l = node638_r & ~pixel[382];
      node695_r = node694_l & pixel[174];
      node695_l = node694_l & ~pixel[174];
      node696_r = node695_l & pixel[377];
      node696_l = node695_l & ~pixel[377];
      node697_r = node696_l & pixel[459];
      node697_l = node696_l & ~pixel[459];
      node698_r = node697_l & pixel[682];
      node698_l = node697_l & ~pixel[682];
      node699 = node698_l;
      node700 = node698_r;
      node701_r = node697_r & pixel[264];
      node701_l = node697_r & ~pixel[264];
      node702 = node701_l;
      node703 = node701_r;
      node704_r = node696_r & pixel[317];
      node704_l = node696_r & ~pixel[317];
      node705_r = node704_l & pixel[633];
      node705_l = node704_l & ~pixel[633];
      node706 = node705_l;
      node707 = node705_r;
      node708_r = node704_r & pixel[556];
      node708_l = node704_r & ~pixel[556];
      node709 = node708_l;
      node710 = node708_r;
      node711_r = node695_r & pixel[268];
      node711_l = node695_r & ~pixel[268];
      node712_r = node711_l & pixel[316];
      node712_l = node711_l & ~pixel[316];
      node713_r = node712_l & pixel[400];
      node713_l = node712_l & ~pixel[400];
      node714 = node713_l;
      node715 = node713_r;
      node716_r = node712_r & pixel[287];
      node716_l = node712_r & ~pixel[287];
      node717 = node716_l;
      node718 = node716_r;
      node719_r = node711_r & pixel[509];
      node719_l = node711_r & ~pixel[509];
      node720 = node719_l;
      node721 = node719_r;
      node722_r = node694_r & pixel[516];
      node722_l = node694_r & ~pixel[516];
      node723_r = node722_l & pixel[464];
      node723_l = node722_l & ~pixel[464];
      node724_r = node723_l & pixel[489];
      node724_l = node723_l & ~pixel[489];
      node725_r = node724_l & pixel[458];
      node725_l = node724_l & ~pixel[458];
      node726 = node725_l;
      node727 = node725_r;
      node728 = node724_r;
      node729_r = node723_r & pixel[567];
      node729_l = node723_r & ~pixel[567];
      node730_r = node729_l & pixel[712];
      node730_l = node729_l & ~pixel[712];
      node731 = node730_l;
      node732 = node730_r;
      node733_r = node729_r & pixel[262];
      node733_l = node729_r & ~pixel[262];
      node734 = node733_l;
      node735 = node733_r;
      node736_r = node722_r & pixel[655];
      node736_l = node722_r & ~pixel[655];
      node737_r = node736_l & pixel[268];
      node737_l = node736_l & ~pixel[268];
      node738_r = node737_l & pixel[244];
      node738_l = node737_l & ~pixel[244];
      node739 = node738_l;
      node740 = node738_r;
      node741_r = node737_r & pixel[660];
      node741_l = node737_r & ~pixel[660];
      node742 = node741_l;
      node743 = node741_r;
      node744_r = node736_r & pixel[175];
      node744_l = node736_r & ~pixel[175];
      node745_r = node744_l & pixel[186];
      node745_l = node744_l & ~pixel[186];
      node746 = node745_l;
      node747 = node745_r;
      node748_r = node744_r & pixel[706];
      node748_l = node744_r & ~pixel[706];
      node749 = node748_l;
      node750 = node748_r;
      node751_r = node637_r & pixel[463];
      node751_l = node637_r & ~pixel[463];
      node752_r = node751_l & pixel[292];
      node752_l = node751_l & ~pixel[292];
      node753_r = node752_l & pixel[191];
      node753_l = node752_l & ~pixel[191];
      node754_r = node753_l & pixel[298];
      node754_l = node753_l & ~pixel[298];
      node755_r = node754_l & pixel[315];
      node755_l = node754_l & ~pixel[315];
      node756_r = node755_l & pixel[345];
      node756_l = node755_l & ~pixel[345];
      node757 = node756_l;
      node758 = node756_r;
      node759_r = node755_r & pixel[178];
      node759_l = node755_r & ~pixel[178];
      node760 = node759_l;
      node761 = node759_r;
      node762_r = node754_r & pixel[653];
      node762_l = node754_r & ~pixel[653];
      node763_r = node762_l & pixel[487];
      node763_l = node762_l & ~pixel[487];
      node764 = node763_l;
      node765 = node763_r;
      node766_r = node762_r & pixel[290];
      node766_l = node762_r & ~pixel[290];
      node767 = node766_l;
      node768 = node766_r;
      node769_r = node753_r & pixel[300];
      node769_l = node753_r & ~pixel[300];
      node770 = node769_l;
      node771_r = node769_r & pixel[633];
      node771_l = node769_r & ~pixel[633];
      node772 = node771_l;
      node773_r = node771_r & pixel[621];
      node773_l = node771_r & ~pixel[621];
      node774 = node773_l;
      node775 = node773_r;
      node776_r = node752_r & pixel[262];
      node776_l = node752_r & ~pixel[262];
      node777_r = node776_l & pixel[150];
      node777_l = node776_l & ~pixel[150];
      node778_r = node777_l & pixel[295];
      node778_l = node777_l & ~pixel[295];
      node779_r = node778_l & pixel[160];
      node779_l = node778_l & ~pixel[160];
      node780 = node779_l;
      node781 = node779_r;
      node782_r = node778_r & pixel[487];
      node782_l = node778_r & ~pixel[487];
      node783 = node782_l;
      node784 = node782_r;
      node785_r = node777_r & pixel[611];
      node785_l = node777_r & ~pixel[611];
      node786_r = node785_l & pixel[261];
      node786_l = node785_l & ~pixel[261];
      node787 = node786_l;
      node788 = node786_r;
      node789 = node785_r;
      node790_r = node776_r & pixel[404];
      node790_l = node776_r & ~pixel[404];
      node791_r = node790_l & pixel[177];
      node791_l = node790_l & ~pixel[177];
      node792_r = node791_l & pixel[242];
      node792_l = node791_l & ~pixel[242];
      node793 = node792_l;
      node794 = node792_r;
      node795_r = node791_r & pixel[461];
      node795_l = node791_r & ~pixel[461];
      node796 = node795_l;
      node797 = node795_r;
      node798_r = node790_r & pixel[432];
      node798_l = node790_r & ~pixel[432];
      node799_r = node798_l & pixel[269];
      node799_l = node798_l & ~pixel[269];
      node800 = node799_l;
      node801 = node799_r;
      node802_r = node798_r & pixel[297];
      node802_l = node798_r & ~pixel[297];
      node803 = node802_l;
      node804 = node802_r;
      node805_r = node751_r & pixel[347];
      node805_l = node751_r & ~pixel[347];
      node806_r = node805_l & pixel[489];
      node806_l = node805_l & ~pixel[489];
      node807_r = node806_l & pixel[628];
      node807_l = node806_l & ~pixel[628];
      node808_r = node807_l & pixel[580];
      node808_l = node807_l & ~pixel[580];
      node809_r = node808_l & pixel[267];
      node809_l = node808_l & ~pixel[267];
      node810 = node809_l;
      node811 = node809_r;
      node812_r = node808_r & pixel[205];
      node812_l = node808_r & ~pixel[205];
      node813 = node812_l;
      node814 = node812_r;
      node815_r = node807_r & pixel[596];
      node815_l = node807_r & ~pixel[596];
      node816_r = node815_l & pixel[405];
      node816_l = node815_l & ~pixel[405];
      node817 = node816_l;
      node818 = node816_r;
      node819_r = node815_r & pixel[523];
      node819_l = node815_r & ~pixel[523];
      node820 = node819_l;
      node821 = node819_r;
      node822_r = node806_r & pixel[154];
      node822_l = node806_r & ~pixel[154];
      node823_r = node822_l & pixel[579];
      node823_l = node822_l & ~pixel[579];
      node824_r = node823_l & pixel[527];
      node824_l = node823_l & ~pixel[527];
      node825 = node824_l;
      node826 = node824_r;
      node827_r = node823_r & pixel[287];
      node827_l = node823_r & ~pixel[287];
      node828 = node827_l;
      node829 = node827_r;
      node830_r = node822_r & pixel[514];
      node830_l = node822_r & ~pixel[514];
      node831_r = node830_l & pixel[516];
      node831_l = node830_l & ~pixel[516];
      node832 = node831_l;
      node833 = node831_r;
      node834_r = node830_r & pixel[349];
      node834_l = node830_r & ~pixel[349];
      node835 = node834_l;
      node836 = node834_r;
      node837_r = node805_r & pixel[487];
      node837_l = node805_r & ~pixel[487];
      node838_r = node837_l & pixel[289];
      node838_l = node837_l & ~pixel[289];
      node839_r = node838_l & pixel[322];
      node839_l = node838_l & ~pixel[322];
      node840_r = node839_l & pixel[579];
      node840_l = node839_l & ~pixel[579];
      node841 = node840_l;
      node842 = node840_r;
      node843_r = node839_r & pixel[517];
      node843_l = node839_r & ~pixel[517];
      node844 = node843_l;
      node845 = node843_r;
      node846_r = node838_r & pixel[516];
      node846_l = node838_r & ~pixel[516];
      node847_r = node846_l & pixel[354];
      node847_l = node846_l & ~pixel[354];
      node848 = node847_l;
      node849 = node847_r;
      node850_r = node846_r & pixel[540];
      node850_l = node846_r & ~pixel[540];
      node851 = node850_l;
      node852 = node850_r;
      node853_r = node837_r & pixel[288];
      node853_l = node837_r & ~pixel[288];
      node854_r = node853_l & pixel[570];
      node854_l = node853_l & ~pixel[570];
      node855_r = node854_l & pixel[185];
      node855_l = node854_l & ~pixel[185];
      node856 = node855_l;
      node857 = node855_r;
      node858_r = node854_r & pixel[460];
      node858_l = node854_r & ~pixel[460];
      node859 = node858_l;
      node860 = node858_r;
      node861_r = node853_r & pixel[96];
      node861_l = node853_r & ~pixel[96];
      node862_r = node861_l & pixel[545];
      node862_l = node861_l & ~pixel[545];
      node863 = node862_l;
      node864 = node862_r;
      node865 = node861_r;
      node866_r = node0_r & pixel[598];
      node866_l = node0_r & ~pixel[598];
      node867_r = node866_l & pixel[69];
      node867_l = node866_l & ~pixel[69];
      node868_r = node867_l & pixel[538];
      node868_l = node867_l & ~pixel[538];
      node869_r = node868_l & pixel[183];
      node869_l = node868_l & ~pixel[183];
      node870_r = node869_l & pixel[570];
      node870_l = node869_l & ~pixel[570];
      node871_r = node870_l & pixel[267];
      node871_l = node870_l & ~pixel[267];
      node872_r = node871_l & pixel[526];
      node872_l = node871_l & ~pixel[526];
      node873_r = node872_l & pixel[571];
      node873_l = node872_l & ~pixel[571];
      node874_r = node873_l & pixel[740];
      node874_l = node873_l & ~pixel[740];
      node875 = node874_l;
      node876 = node874_r;
      node877_r = node873_r & pixel[217];
      node877_l = node873_r & ~pixel[217];
      node878 = node877_l;
      node879 = node877_r;
      node880_r = node872_r & pixel[271];
      node880_l = node872_r & ~pixel[271];
      node881_r = node880_l & pixel[577];
      node881_l = node880_l & ~pixel[577];
      node882 = node881_l;
      node883 = node881_r;
      node884_r = node880_r & pixel[411];
      node884_l = node880_r & ~pixel[411];
      node885 = node884_l;
      node886 = node884_r;
      node887_r = node871_r & pixel[238];
      node887_l = node871_r & ~pixel[238];
      node888_r = node887_l & pixel[430];
      node888_l = node887_l & ~pixel[430];
      node889_r = node888_l & pixel[326];
      node889_l = node888_l & ~pixel[326];
      node890 = node889_l;
      node891 = node889_r;
      node892_r = node888_r & pixel[381];
      node892_l = node888_r & ~pixel[381];
      node893 = node892_l;
      node894 = node892_r;
      node895_r = node887_r & pixel[406];
      node895_l = node887_r & ~pixel[406];
      node896_r = node895_l & pixel[219];
      node896_l = node895_l & ~pixel[219];
      node897 = node896_l;
      node898 = node896_r;
      node899_r = node895_r & pixel[409];
      node899_l = node895_r & ~pixel[409];
      node900 = node899_l;
      node901 = node899_r;
      node902_r = node870_r & pixel[243];
      node902_l = node870_r & ~pixel[243];
      node903_r = node902_l & pixel[241];
      node903_l = node902_l & ~pixel[241];
      node904_r = node903_l & pixel[240];
      node904_l = node903_l & ~pixel[240];
      node905_r = node904_l & pixel[575];
      node905_l = node904_l & ~pixel[575];
      node906 = node905_l;
      node907 = node905_r;
      node908_r = node904_r & pixel[217];
      node908_l = node904_r & ~pixel[217];
      node909 = node908_l;
      node910 = node908_r;
      node911_r = node903_r & pixel[44];
      node911_l = node903_r & ~pixel[44];
      node912_r = node911_l & pixel[657];
      node912_l = node911_l & ~pixel[657];
      node913 = node912_l;
      node914 = node912_r;
      node915_r = node911_r & pixel[264];
      node915_l = node911_r & ~pixel[264];
      node916 = node915_l;
      node917 = node915_r;
      node918_r = node902_r & pixel[180];
      node918_l = node902_r & ~pixel[180];
      node919_r = node918_l & pixel[636];
      node919_l = node918_l & ~pixel[636];
      node920_r = node919_l & pixel[218];
      node920_l = node919_l & ~pixel[218];
      node921 = node920_l;
      node922 = node920_r;
      node923_r = node919_r & pixel[122];
      node923_l = node919_r & ~pixel[122];
      node924 = node923_l;
      node925 = node923_r;
      node926_r = node918_r & pixel[437];
      node926_l = node918_r & ~pixel[437];
      node927_r = node926_l & pixel[348];
      node927_l = node926_l & ~pixel[348];
      node928 = node927_l;
      node929 = node927_r;
      node930 = node926_r;
      node931_r = node869_r & pixel[571];
      node931_l = node869_r & ~pixel[571];
      node932_r = node931_l & pixel[652];
      node932_l = node931_l & ~pixel[652];
      node933_r = node932_l & pixel[581];
      node933_l = node932_l & ~pixel[581];
      node934_r = node933_l & pixel[210];
      node934_l = node933_l & ~pixel[210];
      node935_r = node934_l & pixel[268];
      node935_l = node934_l & ~pixel[268];
      node936 = node935_l;
      node937 = node935_r;
      node938_r = node934_r & pixel[354];
      node938_l = node934_r & ~pixel[354];
      node939 = node938_l;
      node940 = node938_r;
      node941_r = node933_r & pixel[355];
      node941_l = node933_r & ~pixel[355];
      node942_r = node941_l & pixel[351];
      node942_l = node941_l & ~pixel[351];
      node943 = node942_l;
      node944 = node942_r;
      node945_r = node941_r & pixel[632];
      node945_l = node941_r & ~pixel[632];
      node946 = node945_l;
      node947 = node945_r;
      node948_r = node932_r & pixel[379];
      node948_l = node932_r & ~pixel[379];
      node949_r = node948_l & pixel[356];
      node949_l = node948_l & ~pixel[356];
      node950_r = node949_l & pixel[297];
      node950_l = node949_l & ~pixel[297];
      node951 = node950_l;
      node952 = node950_r;
      node953_r = node949_r & pixel[484];
      node953_l = node949_r & ~pixel[484];
      node954 = node953_l;
      node955 = node953_r;
      node956_r = node948_r & pixel[489];
      node956_l = node948_r & ~pixel[489];
      node957_r = node956_l & pixel[345];
      node957_l = node956_l & ~pixel[345];
      node958 = node957_l;
      node959 = node957_r;
      node960_r = node956_r & pixel[678];
      node960_l = node956_r & ~pixel[678];
      node961 = node960_l;
      node962 = node960_r;
      node963_r = node931_r & pixel[299];
      node963_l = node931_r & ~pixel[299];
      node964_r = node963_l & pixel[149];
      node964_l = node963_l & ~pixel[149];
      node965_r = node964_l & pixel[686];
      node965_l = node964_l & ~pixel[686];
      node966_r = node965_l & pixel[297];
      node966_l = node965_l & ~pixel[297];
      node967 = node966_l;
      node968 = node966_r;
      node969_r = node965_r & pixel[516];
      node969_l = node965_r & ~pixel[516];
      node970 = node969_l;
      node971 = node969_r;
      node972_r = node964_r & pixel[438];
      node972_l = node964_r & ~pixel[438];
      node973_r = node972_l & pixel[185];
      node973_l = node972_l & ~pixel[185];
      node974 = node973_l;
      node975 = node973_r;
      node976_r = node972_r & pixel[548];
      node976_l = node972_r & ~pixel[548];
      node977 = node976_l;
      node978 = node976_r;
      node979_r = node963_r & pixel[155];
      node979_l = node963_r & ~pixel[155];
      node980_r = node979_l & pixel[184];
      node980_l = node979_l & ~pixel[184];
      node981_r = node980_l & pixel[260];
      node981_l = node980_l & ~pixel[260];
      node982 = node981_l;
      node983 = node981_r;
      node984_r = node980_r & pixel[496];
      node984_l = node980_r & ~pixel[496];
      node985 = node984_l;
      node986 = node984_r;
      node987_r = node979_r & pixel[213];
      node987_l = node979_r & ~pixel[213];
      node988_r = node987_l & pixel[154];
      node988_l = node987_l & ~pixel[154];
      node989 = node988_l;
      node990 = node988_r;
      node991_r = node987_r & pixel[234];
      node991_l = node987_r & ~pixel[234];
      node992 = node991_l;
      node993 = node991_r;
      node994_r = node868_r & pixel[408];
      node994_l = node868_r & ~pixel[408];
      node995_r = node994_l & pixel[405];
      node995_l = node994_l & ~pixel[405];
      node996_r = node995_l & pixel[487];
      node996_l = node995_l & ~pixel[487];
      node997_r = node996_l & pixel[324];
      node997_l = node996_l & ~pixel[324];
      node998_r = node997_l & pixel[431];
      node998_l = node997_l & ~pixel[431];
      node999_r = node998_l & pixel[566];
      node999_l = node998_l & ~pixel[566];
      node1000 = node999_l;
      node1001 = node999_r;
      node1002_r = node998_r & pixel[434];
      node1002_l = node998_r & ~pixel[434];
      node1003 = node1002_l;
      node1004 = node1002_r;
      node1005_r = node997_r & pixel[455];
      node1005_l = node997_r & ~pixel[455];
      node1006_r = node1005_l & pixel[127];
      node1006_l = node1005_l & ~pixel[127];
      node1007 = node1006_l;
      node1008 = node1006_r;
      node1009_r = node1005_r & pixel[347];
      node1009_l = node1005_r & ~pixel[347];
      node1010 = node1009_l;
      node1011 = node1009_r;
      node1012_r = node996_r & pixel[359];
      node1012_l = node996_r & ~pixel[359];
      node1013_r = node1012_l & pixel[493];
      node1013_l = node1012_l & ~pixel[493];
      node1014_r = node1013_l & pixel[411];
      node1014_l = node1013_l & ~pixel[411];
      node1015 = node1014_l;
      node1016 = node1014_r;
      node1017_r = node1013_r & pixel[156];
      node1017_l = node1013_r & ~pixel[156];
      node1018 = node1017_l;
      node1019 = node1017_r;
      node1020_r = node1012_r & pixel[218];
      node1020_l = node1012_r & ~pixel[218];
      node1021 = node1020_l;
      node1022_r = node1020_r & pixel[627];
      node1022_l = node1020_r & ~pixel[627];
      node1023 = node1022_l;
      node1024 = node1022_r;
      node1025_r = node995_r & pixel[625];
      node1025_l = node995_r & ~pixel[625];
      node1026_r = node1025_l & pixel[248];
      node1026_l = node1025_l & ~pixel[248];
      node1027_r = node1026_l & pixel[183];
      node1027_l = node1026_l & ~pixel[183];
      node1028_r = node1027_l & pixel[455];
      node1028_l = node1027_l & ~pixel[455];
      node1029 = node1028_l;
      node1030 = node1028_r;
      node1031_r = node1027_r & pixel[346];
      node1031_l = node1027_r & ~pixel[346];
      node1032 = node1031_l;
      node1033 = node1031_r;
      node1034_r = node1026_r & pixel[457];
      node1034_l = node1026_r & ~pixel[457];
      node1035 = node1034_l;
      node1036_r = node1034_r & pixel[461];
      node1036_l = node1034_r & ~pixel[461];
      node1037 = node1036_l;
      node1038 = node1036_r;
      node1039_r = node1025_r & pixel[518];
      node1039_l = node1025_r & ~pixel[518];
      node1040_r = node1039_l & pixel[192];
      node1040_l = node1039_l & ~pixel[192];
      node1041_r = node1040_l & pixel[293];
      node1041_l = node1040_l & ~pixel[293];
      node1042 = node1041_l;
      node1043 = node1041_r;
      node1044 = node1040_r;
      node1045_r = node1039_r & pixel[155];
      node1045_l = node1039_r & ~pixel[155];
      node1046_r = node1045_l & pixel[249];
      node1046_l = node1045_l & ~pixel[249];
      node1047 = node1046_l;
      node1048 = node1046_r;
      node1049_r = node1045_r & pixel[457];
      node1049_l = node1045_r & ~pixel[457];
      node1050 = node1049_l;
      node1051 = node1049_r;
      node1052_r = node994_r & pixel[374];
      node1052_l = node994_r & ~pixel[374];
      node1053_r = node1052_l & pixel[341];
      node1053_l = node1052_l & ~pixel[341];
      node1054_r = node1053_l & pixel[650];
      node1054_l = node1053_l & ~pixel[650];
      node1055_r = node1054_l & pixel[652];
      node1055_l = node1054_l & ~pixel[652];
      node1056_r = node1055_l & pixel[370];
      node1056_l = node1055_l & ~pixel[370];
      node1057 = node1056_l;
      node1058 = node1056_r;
      node1059_r = node1055_r & pixel[126];
      node1059_l = node1055_r & ~pixel[126];
      node1060 = node1059_l;
      node1061 = node1059_r;
      node1062_r = node1054_r & pixel[319];
      node1062_l = node1054_r & ~pixel[319];
      node1063_r = node1062_l & pixel[379];
      node1063_l = node1062_l & ~pixel[379];
      node1064 = node1063_l;
      node1065 = node1063_r;
      node1066_r = node1062_r & pixel[348];
      node1066_l = node1062_r & ~pixel[348];
      node1067 = node1066_l;
      node1068 = node1066_r;
      node1069_r = node1053_r & pixel[401];
      node1069_l = node1053_r & ~pixel[401];
      node1070 = node1069_l;
      node1071 = node1069_r;
      node1072_r = node1052_r & pixel[510];
      node1072_l = node1052_r & ~pixel[510];
      node1073_r = node1072_l & pixel[487];
      node1073_l = node1072_l & ~pixel[487];
      node1074_r = node1073_l & pixel[270];
      node1074_l = node1073_l & ~pixel[270];
      node1075_r = node1074_l & pixel[275];
      node1075_l = node1074_l & ~pixel[275];
      node1076 = node1075_l;
      node1077 = node1075_r;
      node1078_r = node1074_r & pixel[343];
      node1078_l = node1074_r & ~pixel[343];
      node1079 = node1078_l;
      node1080 = node1078_r;
      node1081_r = node1073_r & pixel[212];
      node1081_l = node1073_r & ~pixel[212];
      node1082_r = node1081_l & pixel[457];
      node1082_l = node1081_l & ~pixel[457];
      node1083 = node1082_l;
      node1084 = node1082_r;
      node1085_r = node1081_r & pixel[523];
      node1085_l = node1081_r & ~pixel[523];
      node1086 = node1085_l;
      node1087 = node1085_r;
      node1088_r = node1072_r & pixel[683];
      node1088_l = node1072_r & ~pixel[683];
      node1089_r = node1088_l & pixel[291];
      node1089_l = node1088_l & ~pixel[291];
      node1090_r = node1089_l & pixel[541];
      node1090_l = node1089_l & ~pixel[541];
      node1091 = node1090_l;
      node1092 = node1090_r;
      node1093_r = node1089_r & pixel[543];
      node1093_l = node1089_r & ~pixel[543];
      node1094 = node1093_l;
      node1095 = node1093_r;
      node1096_r = node1088_r & pixel[185];
      node1096_l = node1088_r & ~pixel[185];
      node1097_r = node1096_l & pixel[379];
      node1097_l = node1096_l & ~pixel[379];
      node1098 = node1097_l;
      node1099 = node1097_r;
      node1100_r = node1096_r & pixel[489];
      node1100_l = node1096_r & ~pixel[489];
      node1101 = node1100_l;
      node1102 = node1100_r;
      node1103_r = node867_r & pixel[576];
      node1103_l = node867_r & ~pixel[576];
      node1104_r = node1103_l & pixel[234];
      node1104_l = node1103_l & ~pixel[234];
      node1105 = node1104_l;
      node1106 = node1104_r;
      node1107_r = node1103_r & pixel[158];
      node1107_l = node1103_r & ~pixel[158];
      node1108_r = node1107_l & pixel[294];
      node1108_l = node1107_l & ~pixel[294];
      node1109_r = node1108_l & pixel[242];
      node1109_l = node1108_l & ~pixel[242];
      node1110 = node1109_l;
      node1111_r = node1109_r & pixel[371];
      node1111_l = node1109_r & ~pixel[371];
      node1112 = node1111_l;
      node1113 = node1111_r;
      node1114_r = node1108_r & pixel[41];
      node1114_l = node1108_r & ~pixel[41];
      node1115_r = node1114_l & pixel[440];
      node1115_l = node1114_l & ~pixel[440];
      node1116_r = node1115_l & pixel[357];
      node1116_l = node1115_l & ~pixel[357];
      node1117 = node1116_l;
      node1118 = node1116_r;
      node1119 = node1115_r;
      node1120 = node1114_r;
      node1121 = node1107_r;
      node1122_r = node866_r & pixel[483];
      node1122_l = node866_r & ~pixel[483];
      node1123_r = node1122_l & pixel[485];
      node1123_l = node1122_l & ~pixel[485];
      node1124_r = node1123_l & pixel[354];
      node1124_l = node1123_l & ~pixel[354];
      node1125_r = node1124_l & pixel[176];
      node1125_l = node1124_l & ~pixel[176];
      node1126_r = node1125_l & pixel[191];
      node1126_l = node1125_l & ~pixel[191];
      node1127_r = node1126_l & pixel[353];
      node1127_l = node1126_l & ~pixel[353];
      node1128_r = node1127_l & pixel[101];
      node1128_l = node1127_l & ~pixel[101];
      node1129_r = node1128_l & pixel[247];
      node1129_l = node1128_l & ~pixel[247];
      node1130 = node1129_l;
      node1131 = node1129_r;
      node1132_r = node1128_r & pixel[330];
      node1132_l = node1128_r & ~pixel[330];
      node1133 = node1132_l;
      node1134 = node1132_r;
      node1135_r = node1127_r & pixel[263];
      node1135_l = node1127_r & ~pixel[263];
      node1136_r = node1135_l & pixel[350];
      node1136_l = node1135_l & ~pixel[350];
      node1137 = node1136_l;
      node1138 = node1136_r;
      node1139_r = node1135_r & pixel[517];
      node1139_l = node1135_r & ~pixel[517];
      node1140 = node1139_l;
      node1141 = node1139_r;
      node1142_r = node1126_r & pixel[374];
      node1142_l = node1126_r & ~pixel[374];
      node1143_r = node1142_l & pixel[379];
      node1143_l = node1142_l & ~pixel[379];
      node1144_r = node1143_l & pixel[302];
      node1144_l = node1143_l & ~pixel[302];
      node1145 = node1144_l;
      node1146 = node1144_r;
      node1147_r = node1143_r & pixel[489];
      node1147_l = node1143_r & ~pixel[489];
      node1148 = node1147_l;
      node1149 = node1147_r;
      node1150_r = node1142_r & pixel[387];
      node1150_l = node1142_r & ~pixel[387];
      node1151_r = node1150_l & pixel[707];
      node1151_l = node1150_l & ~pixel[707];
      node1152 = node1151_l;
      node1153 = node1151_r;
      node1154 = node1150_r;
      node1155_r = node1125_r & pixel[268];
      node1155_l = node1125_r & ~pixel[268];
      node1156_r = node1155_l & pixel[301];
      node1156_l = node1155_l & ~pixel[301];
      node1157_r = node1156_l & pixel[271];
      node1157_l = node1156_l & ~pixel[271];
      node1158_r = node1157_l & pixel[233];
      node1158_l = node1157_l & ~pixel[233];
      node1159 = node1158_l;
      node1160 = node1158_r;
      node1161_r = node1157_r & pixel[428];
      node1161_l = node1157_r & ~pixel[428];
      node1162 = node1161_l;
      node1163 = node1161_r;
      node1164 = node1156_r;
      node1165_r = node1155_r & pixel[217];
      node1165_l = node1155_r & ~pixel[217];
      node1166_r = node1165_l & pixel[355];
      node1166_l = node1165_l & ~pixel[355];
      node1167_r = node1166_l & pixel[693];
      node1167_l = node1166_l & ~pixel[693];
      node1168 = node1167_l;
      node1169 = node1167_r;
      node1170 = node1166_r;
      node1171_r = node1165_r & pixel[635];
      node1171_l = node1165_r & ~pixel[635];
      node1172_r = node1171_l & pixel[386];
      node1172_l = node1171_l & ~pixel[386];
      node1173 = node1172_l;
      node1174 = node1172_r;
      node1175_r = node1171_r & pixel[235];
      node1175_l = node1171_r & ~pixel[235];
      node1176 = node1175_l;
      node1177 = node1175_r;
      node1178_r = node1124_r & pixel[495];
      node1178_l = node1124_r & ~pixel[495];
      node1179_r = node1178_l & pixel[490];
      node1179_l = node1178_l & ~pixel[490];
      node1180_r = node1179_l & pixel[371];
      node1180_l = node1179_l & ~pixel[371];
      node1181_r = node1180_l & pixel[406];
      node1181_l = node1180_l & ~pixel[406];
      node1182_r = node1181_l & pixel[203];
      node1182_l = node1181_l & ~pixel[203];
      node1183 = node1182_l;
      node1184 = node1182_r;
      node1185_r = node1181_r & pixel[325];
      node1185_l = node1181_r & ~pixel[325];
      node1186 = node1185_l;
      node1187 = node1185_r;
      node1188_r = node1180_r & pixel[658];
      node1188_l = node1180_r & ~pixel[658];
      node1189_r = node1188_l & pixel[238];
      node1189_l = node1188_l & ~pixel[238];
      node1190 = node1189_l;
      node1191 = node1189_r;
      node1192_r = node1188_r & pixel[317];
      node1192_l = node1188_r & ~pixel[317];
      node1193 = node1192_l;
      node1194 = node1192_r;
      node1195_r = node1179_r & pixel[549];
      node1195_l = node1179_r & ~pixel[549];
      node1196_r = node1195_l & pixel[631];
      node1196_l = node1195_l & ~pixel[631];
      node1197_r = node1196_l & pixel[454];
      node1197_l = node1196_l & ~pixel[454];
      node1198 = node1197_l;
      node1199 = node1197_r;
      node1200_r = node1196_r & pixel[472];
      node1200_l = node1196_r & ~pixel[472];
      node1201 = node1200_l;
      node1202 = node1200_r;
      node1203_r = node1195_r & pixel[488];
      node1203_l = node1195_r & ~pixel[488];
      node1204_r = node1203_l & pixel[325];
      node1204_l = node1203_l & ~pixel[325];
      node1205 = node1204_l;
      node1206 = node1204_r;
      node1207_r = node1203_r & pixel[288];
      node1207_l = node1203_r & ~pixel[288];
      node1208 = node1207_l;
      node1209 = node1207_r;
      node1210_r = node1178_r & pixel[318];
      node1210_l = node1178_r & ~pixel[318];
      node1211_r = node1210_l & pixel[629];
      node1211_l = node1210_l & ~pixel[629];
      node1212_r = node1211_l & pixel[454];
      node1212_l = node1211_l & ~pixel[454];
      node1213_r = node1212_l & pixel[591];
      node1213_l = node1212_l & ~pixel[591];
      node1214 = node1213_l;
      node1215 = node1213_r;
      node1216 = node1212_r;
      node1217_r = node1211_r & pixel[377];
      node1217_l = node1211_r & ~pixel[377];
      node1218_r = node1217_l & pixel[400];
      node1218_l = node1217_l & ~pixel[400];
      node1219 = node1218_l;
      node1220 = node1218_r;
      node1221_r = node1217_r & pixel[406];
      node1221_l = node1217_r & ~pixel[406];
      node1222 = node1221_l;
      node1223 = node1221_r;
      node1224_r = node1210_r & pixel[461];
      node1224_l = node1210_r & ~pixel[461];
      node1225_r = node1224_l & pixel[290];
      node1225_l = node1224_l & ~pixel[290];
      node1226_r = node1225_l & pixel[191];
      node1226_l = node1225_l & ~pixel[191];
      node1227 = node1226_l;
      node1228 = node1226_r;
      node1229_r = node1225_r & pixel[346];
      node1229_l = node1225_r & ~pixel[346];
      node1230 = node1229_l;
      node1231 = node1229_r;
      node1232_r = node1224_r & pixel[605];
      node1232_l = node1224_r & ~pixel[605];
      node1233_r = node1232_l & pixel[383];
      node1233_l = node1232_l & ~pixel[383];
      node1234 = node1233_l;
      node1235 = node1233_r;
      node1236_r = node1232_r & pixel[207];
      node1236_l = node1232_r & ~pixel[207];
      node1237 = node1236_l;
      node1238 = node1236_r;
      node1239_r = node1123_r & pixel[655];
      node1239_l = node1123_r & ~pixel[655];
      node1240_r = node1239_l & pixel[548];
      node1240_l = node1239_l & ~pixel[548];
      node1241_r = node1240_l & pixel[623];
      node1241_l = node1240_l & ~pixel[623];
      node1242_r = node1241_l & pixel[659];
      node1242_l = node1241_l & ~pixel[659];
      node1243_r = node1242_l & pixel[604];
      node1243_l = node1242_l & ~pixel[604];
      node1244_r = node1243_l & pixel[290];
      node1244_l = node1243_l & ~pixel[290];
      node1245 = node1244_l;
      node1246 = node1244_r;
      node1247_r = node1243_r & pixel[271];
      node1247_l = node1243_r & ~pixel[271];
      node1248 = node1247_l;
      node1249 = node1247_r;
      node1250_r = node1242_r & pixel[408];
      node1250_l = node1242_r & ~pixel[408];
      node1251_r = node1250_l & pixel[433];
      node1251_l = node1250_l & ~pixel[433];
      node1252 = node1251_l;
      node1253 = node1251_r;
      node1254_r = node1250_r & pixel[235];
      node1254_l = node1250_r & ~pixel[235];
      node1255 = node1254_l;
      node1256 = node1254_r;
      node1257_r = node1241_r & pixel[380];
      node1257_l = node1241_r & ~pixel[380];
      node1258_r = node1257_l & pixel[493];
      node1258_l = node1257_l & ~pixel[493];
      node1259 = node1258_l;
      node1260_r = node1258_r & pixel[381];
      node1260_l = node1258_r & ~pixel[381];
      node1261 = node1260_l;
      node1262 = node1260_r;
      node1263_r = node1257_r & pixel[350];
      node1263_l = node1257_r & ~pixel[350];
      node1264_r = node1263_l & pixel[513];
      node1264_l = node1263_l & ~pixel[513];
      node1265 = node1264_l;
      node1266 = node1264_r;
      node1267_r = node1263_r & pixel[437];
      node1267_l = node1263_r & ~pixel[437];
      node1268 = node1267_l;
      node1269 = node1267_r;
      node1270_r = node1240_r & pixel[216];
      node1270_l = node1240_r & ~pixel[216];
      node1271_r = node1270_l & pixel[612];
      node1271_l = node1270_l & ~pixel[612];
      node1272_r = node1271_l & pixel[241];
      node1272_l = node1271_l & ~pixel[241];
      node1273_r = node1272_l & pixel[473];
      node1273_l = node1272_l & ~pixel[473];
      node1274 = node1273_l;
      node1275 = node1273_r;
      node1276_r = node1272_r & pixel[132];
      node1276_l = node1272_r & ~pixel[132];
      node1277 = node1276_l;
      node1278 = node1276_r;
      node1279 = node1271_r;
      node1280_r = node1270_r & pixel[356];
      node1280_l = node1270_r & ~pixel[356];
      node1281_r = node1280_l & pixel[484];
      node1281_l = node1280_l & ~pixel[484];
      node1282_r = node1281_l & pixel[374];
      node1282_l = node1281_l & ~pixel[374];
      node1283 = node1282_l;
      node1284 = node1282_r;
      node1285_r = node1281_r & pixel[611];
      node1285_l = node1281_r & ~pixel[611];
      node1286 = node1285_l;
      node1287 = node1285_r;
      node1288_r = node1280_r & pixel[426];
      node1288_l = node1280_r & ~pixel[426];
      node1289_r = node1288_l & pixel[407];
      node1289_l = node1288_l & ~pixel[407];
      node1290 = node1289_l;
      node1291 = node1289_r;
      node1292 = node1288_r;
      node1293_r = node1239_r & pixel[324];
      node1293_l = node1239_r & ~pixel[324];
      node1294_r = node1293_l & pixel[299];
      node1294_l = node1293_l & ~pixel[299];
      node1295_r = node1294_l & pixel[329];
      node1295_l = node1294_l & ~pixel[329];
      node1296_r = node1295_l & pixel[570];
      node1296_l = node1295_l & ~pixel[570];
      node1297_r = node1296_l & pixel[544];
      node1297_l = node1296_l & ~pixel[544];
      node1298 = node1297_l;
      node1299 = node1297_r;
      node1300_r = node1296_r & pixel[180];
      node1300_l = node1296_r & ~pixel[180];
      node1301 = node1300_l;
      node1302 = node1300_r;
      node1303_r = node1295_r & pixel[462];
      node1303_l = node1295_r & ~pixel[462];
      node1304_r = node1303_l & pixel[327];
      node1304_l = node1303_l & ~pixel[327];
      node1305 = node1304_l;
      node1306 = node1304_r;
      node1307_r = node1303_r & pixel[456];
      node1307_l = node1303_r & ~pixel[456];
      node1308 = node1307_l;
      node1309 = node1307_r;
      node1310_r = node1294_r & pixel[435];
      node1310_l = node1294_r & ~pixel[435];
      node1311_r = node1310_l & pixel[202];
      node1311_l = node1310_l & ~pixel[202];
      node1312_r = node1311_l & pixel[242];
      node1312_l = node1311_l & ~pixel[242];
      node1313 = node1312_l;
      node1314 = node1312_r;
      node1315 = node1311_r;
      node1316_r = node1310_r & pixel[186];
      node1316_l = node1310_r & ~pixel[186];
      node1317_r = node1316_l & pixel[603];
      node1317_l = node1316_l & ~pixel[603];
      node1318 = node1317_l;
      node1319 = node1317_r;
      node1320_r = node1316_r & pixel[375];
      node1320_l = node1316_r & ~pixel[375];
      node1321 = node1320_l;
      node1322 = node1320_r;
      node1323_r = node1293_r & pixel[432];
      node1323_l = node1293_r & ~pixel[432];
      node1324_r = node1323_l & pixel[268];
      node1324_l = node1323_l & ~pixel[268];
      node1325_r = node1324_l & pixel[487];
      node1325_l = node1324_l & ~pixel[487];
      node1326_r = node1325_l & pixel[316];
      node1326_l = node1325_l & ~pixel[316];
      node1327 = node1326_l;
      node1328 = node1326_r;
      node1329_r = node1325_r & pixel[658];
      node1329_l = node1325_r & ~pixel[658];
      node1330 = node1329_l;
      node1331 = node1329_r;
      node1332_r = node1324_r & pixel[433];
      node1332_l = node1324_r & ~pixel[433];
      node1333_r = node1332_l & pixel[457];
      node1333_l = node1332_l & ~pixel[457];
      node1334 = node1333_l;
      node1335 = node1333_r;
      node1336_r = node1332_r & pixel[548];
      node1336_l = node1332_r & ~pixel[548];
      node1337 = node1336_l;
      node1338 = node1336_r;
      node1339_r = node1323_r & pixel[274];
      node1339_l = node1323_r & ~pixel[274];
      node1340_r = node1339_l & pixel[573];
      node1340_l = node1339_l & ~pixel[573];
      node1341_r = node1340_l & pixel[299];
      node1341_l = node1340_l & ~pixel[299];
      node1342 = node1341_l;
      node1343 = node1341_r;
      node1344_r = node1340_r & pixel[512];
      node1344_l = node1340_r & ~pixel[512];
      node1345 = node1344_l;
      node1346 = node1344_r;
      node1347_r = node1339_r & pixel[592];
      node1347_l = node1339_r & ~pixel[592];
      node1348_r = node1347_l & pixel[541];
      node1348_l = node1347_l & ~pixel[541];
      node1349 = node1348_l;
      node1350 = node1348_r;
      node1351 = node1347_r;
      node1352_r = node1122_r & pixel[318];
      node1352_l = node1122_r & ~pixel[318];
      node1353_r = node1352_l & pixel[267];
      node1353_l = node1352_l & ~pixel[267];
      node1354_r = node1353_l & pixel[655];
      node1354_l = node1353_l & ~pixel[655];
      node1355_r = node1354_l & pixel[214];
      node1355_l = node1354_l & ~pixel[214];
      node1356_r = node1355_l & pixel[442];
      node1356_l = node1355_l & ~pixel[442];
      node1357_r = node1356_l & pixel[158];
      node1357_l = node1356_l & ~pixel[158];
      node1358_r = node1357_l & pixel[124];
      node1358_l = node1357_l & ~pixel[124];
      node1359 = node1358_l;
      node1360 = node1358_r;
      node1361_r = node1357_r & pixel[596];
      node1361_l = node1357_r & ~pixel[596];
      node1362 = node1361_l;
      node1363 = node1361_r;
      node1364_r = node1356_r & pixel[96];
      node1364_l = node1356_r & ~pixel[96];
      node1365_r = node1364_l & pixel[208];
      node1365_l = node1364_l & ~pixel[208];
      node1366 = node1365_l;
      node1367 = node1365_r;
      node1368 = node1364_r;
      node1369_r = node1355_r & pixel[344];
      node1369_l = node1355_r & ~pixel[344];
      node1370_r = node1369_l & pixel[135];
      node1370_l = node1369_l & ~pixel[135];
      node1371_r = node1370_l & pixel[657];
      node1371_l = node1370_l & ~pixel[657];
      node1372 = node1371_l;
      node1373 = node1371_r;
      node1374_r = node1370_r & pixel[347];
      node1374_l = node1370_r & ~pixel[347];
      node1375 = node1374_l;
      node1376 = node1374_r;
      node1377_r = node1369_r & pixel[439];
      node1377_l = node1369_r & ~pixel[439];
      node1378_r = node1377_l & pixel[540];
      node1378_l = node1377_l & ~pixel[540];
      node1379 = node1378_l;
      node1380 = node1378_r;
      node1381_r = node1377_r & pixel[509];
      node1381_l = node1377_r & ~pixel[509];
      node1382 = node1381_l;
      node1383 = node1381_r;
      node1384_r = node1354_r & pixel[624];
      node1384_l = node1354_r & ~pixel[624];
      node1385_r = node1384_l & pixel[379];
      node1385_l = node1384_l & ~pixel[379];
      node1386_r = node1385_l & pixel[409];
      node1386_l = node1385_l & ~pixel[409];
      node1387_r = node1386_l & pixel[200];
      node1387_l = node1386_l & ~pixel[200];
      node1388 = node1387_l;
      node1389 = node1387_r;
      node1390_r = node1386_r & pixel[182];
      node1390_l = node1386_r & ~pixel[182];
      node1391 = node1390_l;
      node1392 = node1390_r;
      node1393_r = node1385_r & pixel[631];
      node1393_l = node1385_r & ~pixel[631];
      node1394_r = node1393_l & pixel[298];
      node1394_l = node1393_l & ~pixel[298];
      node1395 = node1394_l;
      node1396 = node1394_r;
      node1397_r = node1393_r & pixel[151];
      node1397_l = node1393_r & ~pixel[151];
      node1398 = node1397_l;
      node1399 = node1397_r;
      node1400_r = node1384_r & pixel[350];
      node1400_l = node1384_r & ~pixel[350];
      node1401_r = node1400_l & pixel[459];
      node1401_l = node1400_l & ~pixel[459];
      node1402_r = node1401_l & pixel[409];
      node1402_l = node1401_l & ~pixel[409];
      node1403 = node1402_l;
      node1404 = node1402_r;
      node1405_r = node1401_r & pixel[314];
      node1405_l = node1401_r & ~pixel[314];
      node1406 = node1405_l;
      node1407 = node1405_r;
      node1408_r = node1400_r & pixel[461];
      node1408_l = node1400_r & ~pixel[461];
      node1409_r = node1408_l & pixel[551];
      node1409_l = node1408_l & ~pixel[551];
      node1410 = node1409_l;
      node1411 = node1409_r;
      node1412_r = node1408_r & pixel[233];
      node1412_l = node1408_r & ~pixel[233];
      node1413 = node1412_l;
      node1414 = node1412_r;
      node1415_r = node1353_r & pixel[180];
      node1415_l = node1353_r & ~pixel[180];
      node1416_r = node1415_l & pixel[303];
      node1416_l = node1415_l & ~pixel[303];
      node1417_r = node1416_l & pixel[349];
      node1417_l = node1416_l & ~pixel[349];
      node1418_r = node1417_l & pixel[289];
      node1418_l = node1417_l & ~pixel[289];
      node1419_r = node1418_l & pixel[320];
      node1419_l = node1418_l & ~pixel[320];
      node1420 = node1419_l;
      node1421 = node1419_r;
      node1422_r = node1418_r & pixel[602];
      node1422_l = node1418_r & ~pixel[602];
      node1423 = node1422_l;
      node1424 = node1422_r;
      node1425_r = node1417_r & pixel[625];
      node1425_l = node1417_r & ~pixel[625];
      node1426_r = node1425_l & pixel[271];
      node1426_l = node1425_l & ~pixel[271];
      node1427 = node1426_l;
      node1428 = node1426_r;
      node1429_r = node1425_r & pixel[460];
      node1429_l = node1425_r & ~pixel[460];
      node1430 = node1429_l;
      node1431 = node1429_r;
      node1432_r = node1416_r & pixel[381];
      node1432_l = node1416_r & ~pixel[381];
      node1433_r = node1432_l & pixel[494];
      node1433_l = node1432_l & ~pixel[494];
      node1434_r = node1433_l & pixel[134];
      node1434_l = node1433_l & ~pixel[134];
      node1435 = node1434_l;
      node1436 = node1434_r;
      node1437_r = node1433_r & pixel[610];
      node1437_l = node1433_r & ~pixel[610];
      node1438 = node1437_l;
      node1439 = node1437_r;
      node1440_r = node1432_r & pixel[622];
      node1440_l = node1432_r & ~pixel[622];
      node1441_r = node1440_l & pixel[324];
      node1441_l = node1440_l & ~pixel[324];
      node1442 = node1441_l;
      node1443 = node1441_r;
      node1444_r = node1440_r & pixel[345];
      node1444_l = node1440_r & ~pixel[345];
      node1445 = node1444_l;
      node1446 = node1444_r;
      node1447_r = node1415_r & pixel[344];
      node1447_l = node1415_r & ~pixel[344];
      node1448_r = node1447_l & pixel[680];
      node1448_l = node1447_l & ~pixel[680];
      node1449_r = node1448_l & pixel[542];
      node1449_l = node1448_l & ~pixel[542];
      node1450_r = node1449_l & pixel[496];
      node1450_l = node1449_l & ~pixel[496];
      node1451 = node1450_l;
      node1452 = node1450_r;
      node1453_r = node1449_r & pixel[189];
      node1453_l = node1449_r & ~pixel[189];
      node1454 = node1453_l;
      node1455 = node1453_r;
      node1456_r = node1448_r & pixel[514];
      node1456_l = node1448_r & ~pixel[514];
      node1457 = node1456_l;
      node1458_r = node1456_r & pixel[685];
      node1458_l = node1456_r & ~pixel[685];
      node1459 = node1458_l;
      node1460 = node1458_r;
      node1461_r = node1447_r & pixel[407];
      node1461_l = node1447_r & ~pixel[407];
      node1462_r = node1461_l & pixel[374];
      node1462_l = node1461_l & ~pixel[374];
      node1463 = node1462_l;
      node1464_r = node1462_r & pixel[554];
      node1464_l = node1462_r & ~pixel[554];
      node1465 = node1464_l;
      node1466 = node1464_r;
      node1467_r = node1461_r & pixel[654];
      node1467_l = node1461_r & ~pixel[654];
      node1468_r = node1467_l & pixel[521];
      node1468_l = node1467_l & ~pixel[521];
      node1469 = node1468_l;
      node1470 = node1468_r;
      node1471_r = node1467_r & pixel[454];
      node1471_l = node1467_r & ~pixel[454];
      node1472 = node1471_l;
      node1473 = node1471_r;
      node1474_r = node1352_r & pixel[461];
      node1474_l = node1352_r & ~pixel[461];
      node1475_r = node1474_l & pixel[242];
      node1475_l = node1474_l & ~pixel[242];
      node1476_r = node1475_l & pixel[273];
      node1476_l = node1475_l & ~pixel[273];
      node1477_r = node1476_l & pixel[657];
      node1477_l = node1476_l & ~pixel[657];
      node1478_r = node1477_l & pixel[274];
      node1478_l = node1477_l & ~pixel[274];
      node1479_r = node1478_l & pixel[135];
      node1479_l = node1478_l & ~pixel[135];
      node1480 = node1479_l;
      node1481 = node1479_r;
      node1482_r = node1478_r & pixel[379];
      node1482_l = node1478_r & ~pixel[379];
      node1483 = node1482_l;
      node1484 = node1482_r;
      node1485_r = node1477_r & pixel[409];
      node1485_l = node1477_r & ~pixel[409];
      node1486_r = node1485_l & pixel[372];
      node1486_l = node1485_l & ~pixel[372];
      node1487 = node1486_l;
      node1488 = node1486_r;
      node1489_r = node1485_r & pixel[457];
      node1489_l = node1485_r & ~pixel[457];
      node1490 = node1489_l;
      node1491 = node1489_r;
      node1492_r = node1476_r & pixel[428];
      node1492_l = node1476_r & ~pixel[428];
      node1493_r = node1492_l & pixel[514];
      node1493_l = node1492_l & ~pixel[514];
      node1494_r = node1493_l & pixel[207];
      node1494_l = node1493_l & ~pixel[207];
      node1495 = node1494_l;
      node1496 = node1494_r;
      node1497_r = node1493_r & pixel[247];
      node1497_l = node1493_r & ~pixel[247];
      node1498 = node1497_l;
      node1499 = node1497_r;
      node1500_r = node1492_r & pixel[626];
      node1500_l = node1492_r & ~pixel[626];
      node1501_r = node1500_l & pixel[231];
      node1501_l = node1500_l & ~pixel[231];
      node1502 = node1501_l;
      node1503 = node1501_r;
      node1504_r = node1500_r & pixel[357];
      node1504_l = node1500_r & ~pixel[357];
      node1505 = node1504_l;
      node1506 = node1504_r;
      node1507_r = node1475_r & pixel[495];
      node1507_l = node1475_r & ~pixel[495];
      node1508_r = node1507_l & pixel[352];
      node1508_l = node1507_l & ~pixel[352];
      node1509_r = node1508_l & pixel[219];
      node1509_l = node1508_l & ~pixel[219];
      node1510_r = node1509_l & pixel[488];
      node1510_l = node1509_l & ~pixel[488];
      node1511 = node1510_l;
      node1512 = node1510_r;
      node1513_r = node1509_r & pixel[359];
      node1513_l = node1509_r & ~pixel[359];
      node1514 = node1513_l;
      node1515 = node1513_r;
      node1516_r = node1508_r & pixel[378];
      node1516_l = node1508_r & ~pixel[378];
      node1517_r = node1516_l & pixel[369];
      node1517_l = node1516_l & ~pixel[369];
      node1518 = node1517_l;
      node1519 = node1517_r;
      node1520_r = node1516_r & pixel[274];
      node1520_l = node1516_r & ~pixel[274];
      node1521 = node1520_l;
      node1522 = node1520_r;
      node1523_r = node1507_r & pixel[713];
      node1523_l = node1507_r & ~pixel[713];
      node1524_r = node1523_l & pixel[428];
      node1524_l = node1523_l & ~pixel[428];
      node1525_r = node1524_l & pixel[415];
      node1525_l = node1524_l & ~pixel[415];
      node1526 = node1525_l;
      node1527 = node1525_r;
      node1528_r = node1524_r & pixel[173];
      node1528_l = node1524_r & ~pixel[173];
      node1529 = node1528_l;
      node1530 = node1528_r;
      node1531_r = node1523_r & pixel[443];
      node1531_l = node1523_r & ~pixel[443];
      node1532 = node1531_l;
      node1533 = node1531_r;
      node1534_r = node1474_r & pixel[549];
      node1534_l = node1474_r & ~pixel[549];
      node1535_r = node1534_l & pixel[399];
      node1535_l = node1534_l & ~pixel[399];
      node1536_r = node1535_l & pixel[184];
      node1536_l = node1535_l & ~pixel[184];
      node1537_r = node1536_l & pixel[427];
      node1537_l = node1536_l & ~pixel[427];
      node1538_r = node1537_l & pixel[412];
      node1538_l = node1537_l & ~pixel[412];
      node1539 = node1538_l;
      node1540 = node1538_r;
      node1541_r = node1537_r & pixel[162];
      node1541_l = node1537_r & ~pixel[162];
      node1542 = node1541_l;
      node1543 = node1541_r;
      node1544_r = node1536_r & pixel[131];
      node1544_l = node1536_r & ~pixel[131];
      node1545_r = node1544_l & pixel[521];
      node1545_l = node1544_l & ~pixel[521];
      node1546 = node1545_l;
      node1547 = node1545_r;
      node1548_r = node1544_r & pixel[624];
      node1548_l = node1544_r & ~pixel[624];
      node1549 = node1548_l;
      node1550 = node1548_r;
      node1551_r = node1535_r & pixel[580];
      node1551_l = node1535_r & ~pixel[580];
      node1552_r = node1551_l & pixel[737];
      node1552_l = node1551_l & ~pixel[737];
      node1553_r = node1552_l & pixel[239];
      node1553_l = node1552_l & ~pixel[239];
      node1554 = node1553_l;
      node1555 = node1553_r;
      node1556 = node1552_r;
      node1557_r = node1551_r & pixel[595];
      node1557_l = node1551_r & ~pixel[595];
      node1558 = node1557_l;
      node1559_r = node1557_r & pixel[260];
      node1559_l = node1557_r & ~pixel[260];
      node1560 = node1559_l;
      node1561 = node1559_r;
      node1562_r = node1534_r & pixel[655];
      node1562_l = node1534_r & ~pixel[655];
      node1563_r = node1562_l & pixel[219];
      node1563_l = node1562_l & ~pixel[219];
      node1564_r = node1563_l & pixel[245];
      node1564_l = node1563_l & ~pixel[245];
      node1565_r = node1564_l & pixel[611];
      node1565_l = node1564_l & ~pixel[611];
      node1566 = node1565_l;
      node1567 = node1565_r;
      node1568_r = node1564_r & pixel[150];
      node1568_l = node1564_r & ~pixel[150];
      node1569 = node1568_l;
      node1570 = node1568_r;
      node1571_r = node1563_r & pixel[453];
      node1571_l = node1563_r & ~pixel[453];
      node1572_r = node1571_l & pixel[125];
      node1572_l = node1571_l & ~pixel[125];
      node1573 = node1572_l;
      node1574 = node1572_r;
      node1575_r = node1571_r & pixel[488];
      node1575_l = node1571_r & ~pixel[488];
      node1576 = node1575_l;
      node1577 = node1575_r;
      node1578_r = node1562_r & pixel[385];
      node1578_l = node1562_r & ~pixel[385];
      node1579_r = node1578_l & pixel[354];
      node1579_l = node1578_l & ~pixel[354];
      node1580_r = node1579_l & pixel[684];
      node1580_l = node1579_l & ~pixel[684];
      node1581 = node1580_l;
      node1582 = node1580_r;
      node1583_r = node1579_r & pixel[426];
      node1583_l = node1579_r & ~pixel[426];
      node1584 = node1583_l;
      node1585 = node1583_r;
      node1586_r = node1578_r & pixel[523];
      node1586_l = node1578_r & ~pixel[523];
      node1587_r = node1586_l & pixel[683];
      node1587_l = node1586_l & ~pixel[683];
      node1588 = node1587_l;
      node1589 = node1587_r;
      node1590_r = node1586_r & pixel[552];
      node1590_l = node1586_r & ~pixel[552];
      node1591 = node1590_l;
      node1592 = node1590_r;
      result0 = node32 | node76 | node81 | node83 | node91 | node102 | node103 | node113 | node143 | node147 | node148 | node236 | node240 | node255 | node267 | node318 | node369 | node372 | node374 | node378 | node400 | node408 | node425 | node451 | node470 | node558 | node572 | node647 | node648 | node682 | node910 | node917 | node921 | node928 | node955 | node1000 | node1001 | node1003 | node1011 | node1021 | node1024 | node1037 | node1043 | node1050 | node1120 | node1249 | node1252 | node1290 | node1305 | node1313 | node1314 | node1331 | node1335 | node1380 | node1382 | node1388 | node1403 | node1430 | node1438 | node1446 | node1459 | node1463 | node1466 | node1469 | node1481 | node1483 | node1488 | node1498 | node1505 | node1506 | node1511 | node1512 | node1515 | node1518 | node1519 | node1522 | node1527 | node1529 | node1533 | node1577 | node1588 | node1591 | node1592;
      result1 = node10 | node17 | node121 | node217 | node224 | node225 | node233 | node247 | node253 | node260 | node287 | node342 | node344 | node391 | node1268 | node1375;
      result2 = node11 | node14 | node20 | node21 | node25 | node28 | node96 | node165 | node228 | node341 | node350 | node357 | node360 | node366 | node388 | node390 | node392 | node396 | node427 | node455 | node456 | node464 | node492 | node500 | node506 | node516 | node520 | node531 | node607 | node616 | node623 | node645 | node671 | node675 | node679 | node681 | node686 | node692 | node702 | node734 | node740 | node742 | node813 | node826 | node835 | node852 | node909 | node916 | node925 | node968 | node974 | node1004 | node1008 | node1010 | node1016 | node1019 | node1030 | node1032 | node1033 | node1042 | node1057 | node1061 | node1064 | node1083 | node1092 | node1105 | node1112 | node1117 | node1121 | node1134 | node1146 | node1154 | node1170 | node1205 | node1216 | node1245 | node1253 | node1275 | node1277 | node1279 | node1287 | node1292 | node1360 | node1362 | node1363 | node1367 | node1372 | node1373 | node1383 | node1389 | node1392 | node1404 | node1406 | node1414 | node1420 | node1421 | node1423 | node1428 | node1452 | node1454 | node1455 | node1470 | node1473 | node1547 | node1550 | node1567 | node1569;
      result3 = node26 | node36 | node45 | node128 | node170 | node172 | node173 | node177 | node218 | node220 | node283 | node295 | node301 | node313 | node319 | node321 | node322 | node327 | node335 | node337 | node338 | node365 | node387 | node397 | node402 | node404 | node421 | node433 | node440 | node449 | node458 | node484 | node486 | node498 | node499 | node508 | node542 | node544 | node554 | node574 | node626 | node666 | node700 | node707 | node714 | node717 | node720 | node735 | node757 | node764 | node767 | node768 | node772 | node775 | node783 | node787 | node788 | node814 | node818 | node820 | node821 | node828 | node832 | node833 | node842 | node844 | node845 | node857 | node944 | node958 | node962 | node1067 | node1079 | node1101 | node1138 | node1148 | node1159 | node1162 | node1168 | node1173 | node1184 | node1186 | node1187 | node1193 | node1206 | node1208 | node1215 | node1219 | node1222 | node1223 | node1227 | node1228 | node1230 | node1238 | node1283 | node1334 | node1342 | node1345 | node1351 | node1399 | node1411 | node1457 | node1496 | node1530;
      result4 = node73 | node77 | node109 | node124 | node179 | node186 | node188 | node424 | node476 | node491 | node521 | node527 | node541 | node546 | node578 | node588 | node595 | node596 | node600 | node631 | node655 | node672 | node690 | node731 | node841 | node875 | node879 | node882 | node885 | node886 | node894 | node924 | node930 | node937 | node982 | node989 | node1018 | node1023 | node1058 | node1071 | node1084 | node1091 | node1094 | node1095 | node1099 | node1137 | node1141 | node1149 | node1199 | node1234 | node1235 | node1246 | node1265 | node1299 | node1318 | node1330 | node1337 | node1349 | node1359 | node1376 | node1391 | node1396 | node1542 | node1543 | node1554 | node1555 | node1585;
      result5 = node41 | node59 | node63 | node66 | node104 | node105 | node122 | node129 | node131 | node139 | node140 | node144 | node146 | node154 | node157 | node161 | node162 | node164 | node232 | node250 | node262 | node266 | node276 | node294 | node302 | node307 | node308 | node324 | node326 | node368 | node405 | node436 | node442 | node448 | node452 | node463 | node469 | node483 | node487 | node523 | node528 | node539 | node547 | node552 | node555 | node589 | node609 | node644 | node699 | node709 | node715 | node718 | node721 | node726 | node758 | node761 | node770 | node780 | node781 | node789 | node793 | node794 | node796 | node800 | node801 | node803 | node848 | node890 | node893 | node898 | node900 | node922 | node943 | node951 | node952 | node959 | node970 | node977 | node1007 | node1015 | node1029 | node1035 | node1044 | node1048 | node1076 | node1130 | node1131 | node1140 | node1145 | node1152 | node1160 | node1163 | node1177 | node1183 | node1194 | node1231 | node1259 | node1284 | node1298 | node1302 | node1306 | node1328 | node1338 | node1395 | node1435 | node1442 | node1465 | node1490 | node1491 | node1514 | node1526 | node1539 | node1573 | node1581 | node1582;
      result6 = node35 | node74 | node84 | node89 | node92 | node95 | node97 | node110 | node114 | node132 | node185 | node198 | node291 | node352 | node353 | node373 | node379 | node381 | node399 | node407 | node479 | node505 | node524 | node559 | node573 | node678 | node703 | node706 | node710 | node739 | node856 | node865 | node878 | node883 | node906 | node907 | node913 | node929 | node967 | node978 | node990 | node1106 | node1110 | node1113 | node1118 | node1119 | node1133 | node1248 | node1255 | node1261 | node1274 | node1278 | node1286 | node1301 | node1366 | node1368 | node1424 | node1427 | node1431 | node1480 | node1502 | node1549 | node1558 | node1560 | node1566 | node1570 | node1574;
      result7 = node13 | node18 | node29 | node48 | node80 | node137 | node193 | node194 | node227 | node241 | node246 | node277 | node279 | node298 | node334 | node380 | node417 | node420 | node435 | node439 | node443 | node465 | node467 | node538 | node551 | node566 | node568 | node569 | node579 | node582 | node585 | node597 | node601 | node606 | node610 | node617 | node622 | node630 | node635 | node651 | node654 | node658 | node661 | node665 | node693 | node750 | node811 | node817 | node825 | node891 | node897 | node983 | node1098 | node1202 | node1214 | node1269 | node1540;
      result8 = node42 | node44 | node56 | node57 | node67 | node112 | node125 | node136 | node158 | node180 | node189 | node192 | node199 | node201 | node202 | node205 | node206 | node208 | node209 | node221 | node235 | node239 | node249 | node254 | node259 | node263 | node269 | node270 | node284 | node286 | node292 | node299 | node310 | node311 | node314 | node345 | node349 | node356 | node359 | node459 | node509 | node512 | node513 | node530 | node634 | node636 | node727 | node728 | node743 | node746 | node747 | node749 | node760 | node765 | node774 | node784 | node797 | node804 | node836 | node851 | node859 | node860 | node863 | node864 | node914 | node947 | node954 | node961 | node971 | node975 | node993 | node1038 | node1047 | node1051 | node1060 | node1065 | node1068 | node1077 | node1086 | node1087 | node1102 | node1174 | node1176 | node1190 | node1201 | node1209 | node1220 | node1237 | node1256 | node1266 | node1291 | node1308 | node1315 | node1319 | node1321 | node1322 | node1327 | node1343 | node1346 | node1350 | node1379 | node1398 | node1410 | node1413 | node1436 | node1439 | node1443 | node1445 | node1451 | node1460 | node1472 | node1484 | node1487 | node1495 | node1499 | node1503 | node1521 | node1532 | node1546 | node1561 | node1576 | node1584 | node1589;
      result9 = node33 | node49 | node51 | node52 | node60 | node64 | node88 | node155 | node169 | node176 | node280 | node418 | node428 | node432 | node477 | node480 | node494 | node495 | node515 | node560 | node565 | node581 | node586 | node602 | node613 | node614 | node625 | node627 | node652 | node660 | node664 | node674 | node687 | node689 | node732 | node810 | node829 | node849 | node876 | node901 | node936 | node939 | node940 | node946 | node985 | node986 | node992 | node1070 | node1080 | node1153 | node1164 | node1169 | node1191 | node1198 | node1262 | node1309 | node1407 | node1556;

      tree_8 = {result9, result8, result7, result6, result5, result4, result3, result2, result1, result0};
    end
  endfunction

  function [9:0] tree_9;
    input [783:0] pixel;

    reg node0_r;
    reg node0_l;
    reg node1_r;
    reg node1_l;
    reg node2_r;
    reg node2_l;
    reg node3_r;
    reg node3_l;
    reg node4_r;
    reg node4_l;
    reg node5_r;
    reg node5_l;
    reg node6_r;
    reg node6_l;
    reg node7_r;
    reg node7_l;
    reg node8_r;
    reg node8_l;
    reg node9_r;
    reg node9_l;
    reg node10;
    reg node11;
    reg node12_r;
    reg node12_l;
    reg node13;
    reg node14;
    reg node15_r;
    reg node15_l;
    reg node16_r;
    reg node16_l;
    reg node17;
    reg node18;
    reg node19_r;
    reg node19_l;
    reg node20;
    reg node21;
    reg node22_r;
    reg node22_l;
    reg node23_r;
    reg node23_l;
    reg node24_r;
    reg node24_l;
    reg node25;
    reg node26;
    reg node27_r;
    reg node27_l;
    reg node28;
    reg node29;
    reg node30_r;
    reg node30_l;
    reg node31_r;
    reg node31_l;
    reg node32;
    reg node33;
    reg node34_r;
    reg node34_l;
    reg node35;
    reg node36;
    reg node37_r;
    reg node37_l;
    reg node38_r;
    reg node38_l;
    reg node39_r;
    reg node39_l;
    reg node40_r;
    reg node40_l;
    reg node41;
    reg node42;
    reg node43_r;
    reg node43_l;
    reg node44;
    reg node45;
    reg node46_r;
    reg node46_l;
    reg node47;
    reg node48_r;
    reg node48_l;
    reg node49;
    reg node50;
    reg node51_r;
    reg node51_l;
    reg node52_r;
    reg node52_l;
    reg node53_r;
    reg node53_l;
    reg node54;
    reg node55;
    reg node56_r;
    reg node56_l;
    reg node57;
    reg node58;
    reg node59_r;
    reg node59_l;
    reg node60;
    reg node61;
    reg node62_r;
    reg node62_l;
    reg node63_r;
    reg node63_l;
    reg node64_r;
    reg node64_l;
    reg node65_r;
    reg node65_l;
    reg node66_r;
    reg node66_l;
    reg node67;
    reg node68;
    reg node69_r;
    reg node69_l;
    reg node70;
    reg node71;
    reg node72_r;
    reg node72_l;
    reg node73_r;
    reg node73_l;
    reg node74;
    reg node75;
    reg node76_r;
    reg node76_l;
    reg node77;
    reg node78;
    reg node79_r;
    reg node79_l;
    reg node80_r;
    reg node80_l;
    reg node81_r;
    reg node81_l;
    reg node82;
    reg node83;
    reg node84_r;
    reg node84_l;
    reg node85;
    reg node86;
    reg node87_r;
    reg node87_l;
    reg node88_r;
    reg node88_l;
    reg node89;
    reg node90;
    reg node91;
    reg node92_r;
    reg node92_l;
    reg node93_r;
    reg node93_l;
    reg node94_r;
    reg node94_l;
    reg node95_r;
    reg node95_l;
    reg node96;
    reg node97;
    reg node98_r;
    reg node98_l;
    reg node99;
    reg node100;
    reg node101_r;
    reg node101_l;
    reg node102_r;
    reg node102_l;
    reg node103;
    reg node104;
    reg node105_r;
    reg node105_l;
    reg node106;
    reg node107;
    reg node108_r;
    reg node108_l;
    reg node109_r;
    reg node109_l;
    reg node110_r;
    reg node110_l;
    reg node111;
    reg node112;
    reg node113_r;
    reg node113_l;
    reg node114;
    reg node115;
    reg node116_r;
    reg node116_l;
    reg node117_r;
    reg node117_l;
    reg node118;
    reg node119;
    reg node120;
    reg node121_r;
    reg node121_l;
    reg node122_r;
    reg node122_l;
    reg node123_r;
    reg node123_l;
    reg node124_r;
    reg node124_l;
    reg node125_r;
    reg node125_l;
    reg node126_r;
    reg node126_l;
    reg node127;
    reg node128;
    reg node129_r;
    reg node129_l;
    reg node130;
    reg node131;
    reg node132_r;
    reg node132_l;
    reg node133_r;
    reg node133_l;
    reg node134;
    reg node135;
    reg node136_r;
    reg node136_l;
    reg node137;
    reg node138;
    reg node139_r;
    reg node139_l;
    reg node140_r;
    reg node140_l;
    reg node141_r;
    reg node141_l;
    reg node142;
    reg node143;
    reg node144_r;
    reg node144_l;
    reg node145;
    reg node146;
    reg node147_r;
    reg node147_l;
    reg node148_r;
    reg node148_l;
    reg node149;
    reg node150;
    reg node151_r;
    reg node151_l;
    reg node152;
    reg node153;
    reg node154_r;
    reg node154_l;
    reg node155_r;
    reg node155_l;
    reg node156;
    reg node157;
    reg node158_r;
    reg node158_l;
    reg node159_r;
    reg node159_l;
    reg node160_r;
    reg node160_l;
    reg node161;
    reg node162;
    reg node163_r;
    reg node163_l;
    reg node164;
    reg node165;
    reg node166_r;
    reg node166_l;
    reg node167;
    reg node168;
    reg node169_r;
    reg node169_l;
    reg node170_r;
    reg node170_l;
    reg node171_r;
    reg node171_l;
    reg node172_r;
    reg node172_l;
    reg node173_r;
    reg node173_l;
    reg node174;
    reg node175;
    reg node176_r;
    reg node176_l;
    reg node177;
    reg node178;
    reg node179;
    reg node180_r;
    reg node180_l;
    reg node181_r;
    reg node181_l;
    reg node182_r;
    reg node182_l;
    reg node183;
    reg node184;
    reg node185_r;
    reg node185_l;
    reg node186;
    reg node187;
    reg node188_r;
    reg node188_l;
    reg node189_r;
    reg node189_l;
    reg node190;
    reg node191;
    reg node192_r;
    reg node192_l;
    reg node193;
    reg node194;
    reg node195_r;
    reg node195_l;
    reg node196_r;
    reg node196_l;
    reg node197;
    reg node198_r;
    reg node198_l;
    reg node199;
    reg node200;
    reg node201;
    reg node202_r;
    reg node202_l;
    reg node203_r;
    reg node203_l;
    reg node204_r;
    reg node204_l;
    reg node205_r;
    reg node205_l;
    reg node206_r;
    reg node206_l;
    reg node207_r;
    reg node207_l;
    reg node208_r;
    reg node208_l;
    reg node209;
    reg node210;
    reg node211_r;
    reg node211_l;
    reg node212;
    reg node213;
    reg node214_r;
    reg node214_l;
    reg node215_r;
    reg node215_l;
    reg node216;
    reg node217;
    reg node218_r;
    reg node218_l;
    reg node219;
    reg node220;
    reg node221_r;
    reg node221_l;
    reg node222_r;
    reg node222_l;
    reg node223_r;
    reg node223_l;
    reg node224;
    reg node225;
    reg node226_r;
    reg node226_l;
    reg node227;
    reg node228;
    reg node229_r;
    reg node229_l;
    reg node230_r;
    reg node230_l;
    reg node231;
    reg node232;
    reg node233;
    reg node234_r;
    reg node234_l;
    reg node235_r;
    reg node235_l;
    reg node236_r;
    reg node236_l;
    reg node237_r;
    reg node237_l;
    reg node238;
    reg node239;
    reg node240_r;
    reg node240_l;
    reg node241;
    reg node242;
    reg node243;
    reg node244_r;
    reg node244_l;
    reg node245_r;
    reg node245_l;
    reg node246_r;
    reg node246_l;
    reg node247;
    reg node248;
    reg node249_r;
    reg node249_l;
    reg node250;
    reg node251;
    reg node252_r;
    reg node252_l;
    reg node253_r;
    reg node253_l;
    reg node254;
    reg node255;
    reg node256_r;
    reg node256_l;
    reg node257;
    reg node258;
    reg node259_r;
    reg node259_l;
    reg node260_r;
    reg node260_l;
    reg node261_r;
    reg node261_l;
    reg node262_r;
    reg node262_l;
    reg node263_r;
    reg node263_l;
    reg node264;
    reg node265;
    reg node266_r;
    reg node266_l;
    reg node267;
    reg node268;
    reg node269_r;
    reg node269_l;
    reg node270_r;
    reg node270_l;
    reg node271;
    reg node272;
    reg node273;
    reg node274_r;
    reg node274_l;
    reg node275_r;
    reg node275_l;
    reg node276_r;
    reg node276_l;
    reg node277;
    reg node278;
    reg node279;
    reg node280_r;
    reg node280_l;
    reg node281;
    reg node282_r;
    reg node282_l;
    reg node283;
    reg node284;
    reg node285_r;
    reg node285_l;
    reg node286_r;
    reg node286_l;
    reg node287_r;
    reg node287_l;
    reg node288_r;
    reg node288_l;
    reg node289;
    reg node290;
    reg node291_r;
    reg node291_l;
    reg node292;
    reg node293;
    reg node294_r;
    reg node294_l;
    reg node295_r;
    reg node295_l;
    reg node296;
    reg node297;
    reg node298_r;
    reg node298_l;
    reg node299;
    reg node300;
    reg node301_r;
    reg node301_l;
    reg node302_r;
    reg node302_l;
    reg node303_r;
    reg node303_l;
    reg node304;
    reg node305;
    reg node306;
    reg node307_r;
    reg node307_l;
    reg node308_r;
    reg node308_l;
    reg node309;
    reg node310;
    reg node311_r;
    reg node311_l;
    reg node312;
    reg node313;
    reg node314_r;
    reg node314_l;
    reg node315_r;
    reg node315_l;
    reg node316_r;
    reg node316_l;
    reg node317_r;
    reg node317_l;
    reg node318_r;
    reg node318_l;
    reg node319_r;
    reg node319_l;
    reg node320;
    reg node321;
    reg node322_r;
    reg node322_l;
    reg node323;
    reg node324;
    reg node325_r;
    reg node325_l;
    reg node326_r;
    reg node326_l;
    reg node327;
    reg node328;
    reg node329_r;
    reg node329_l;
    reg node330;
    reg node331;
    reg node332;
    reg node333_r;
    reg node333_l;
    reg node334_r;
    reg node334_l;
    reg node335_r;
    reg node335_l;
    reg node336_r;
    reg node336_l;
    reg node337;
    reg node338;
    reg node339_r;
    reg node339_l;
    reg node340;
    reg node341;
    reg node342_r;
    reg node342_l;
    reg node343;
    reg node344_r;
    reg node344_l;
    reg node345;
    reg node346;
    reg node347_r;
    reg node347_l;
    reg node348_r;
    reg node348_l;
    reg node349_r;
    reg node349_l;
    reg node350;
    reg node351;
    reg node352_r;
    reg node352_l;
    reg node353;
    reg node354;
    reg node355_r;
    reg node355_l;
    reg node356;
    reg node357_r;
    reg node357_l;
    reg node358;
    reg node359;
    reg node360_r;
    reg node360_l;
    reg node361_r;
    reg node361_l;
    reg node362_r;
    reg node362_l;
    reg node363_r;
    reg node363_l;
    reg node364_r;
    reg node364_l;
    reg node365;
    reg node366;
    reg node367_r;
    reg node367_l;
    reg node368;
    reg node369;
    reg node370_r;
    reg node370_l;
    reg node371_r;
    reg node371_l;
    reg node372;
    reg node373;
    reg node374;
    reg node375_r;
    reg node375_l;
    reg node376_r;
    reg node376_l;
    reg node377_r;
    reg node377_l;
    reg node378;
    reg node379;
    reg node380_r;
    reg node380_l;
    reg node381;
    reg node382;
    reg node383_r;
    reg node383_l;
    reg node384_r;
    reg node384_l;
    reg node385;
    reg node386;
    reg node387_r;
    reg node387_l;
    reg node388;
    reg node389;
    reg node390_r;
    reg node390_l;
    reg node391_r;
    reg node391_l;
    reg node392_r;
    reg node392_l;
    reg node393_r;
    reg node393_l;
    reg node394;
    reg node395;
    reg node396_r;
    reg node396_l;
    reg node397;
    reg node398;
    reg node399_r;
    reg node399_l;
    reg node400_r;
    reg node400_l;
    reg node401;
    reg node402;
    reg node403;
    reg node404_r;
    reg node404_l;
    reg node405_r;
    reg node405_l;
    reg node406;
    reg node407_r;
    reg node407_l;
    reg node408;
    reg node409;
    reg node410_r;
    reg node410_l;
    reg node411;
    reg node412;
    reg node413_r;
    reg node413_l;
    reg node414_r;
    reg node414_l;
    reg node415_r;
    reg node415_l;
    reg node416_r;
    reg node416_l;
    reg node417_r;
    reg node417_l;
    reg node418_r;
    reg node418_l;
    reg node419_r;
    reg node419_l;
    reg node420_r;
    reg node420_l;
    reg node421;
    reg node422;
    reg node423_r;
    reg node423_l;
    reg node424;
    reg node425;
    reg node426_r;
    reg node426_l;
    reg node427_r;
    reg node427_l;
    reg node428;
    reg node429;
    reg node430_r;
    reg node430_l;
    reg node431;
    reg node432;
    reg node433_r;
    reg node433_l;
    reg node434_r;
    reg node434_l;
    reg node435_r;
    reg node435_l;
    reg node436;
    reg node437;
    reg node438_r;
    reg node438_l;
    reg node439;
    reg node440;
    reg node441_r;
    reg node441_l;
    reg node442_r;
    reg node442_l;
    reg node443;
    reg node444;
    reg node445_r;
    reg node445_l;
    reg node446;
    reg node447;
    reg node448_r;
    reg node448_l;
    reg node449_r;
    reg node449_l;
    reg node450_r;
    reg node450_l;
    reg node451_r;
    reg node451_l;
    reg node452;
    reg node453;
    reg node454_r;
    reg node454_l;
    reg node455;
    reg node456;
    reg node457_r;
    reg node457_l;
    reg node458_r;
    reg node458_l;
    reg node459;
    reg node460;
    reg node461_r;
    reg node461_l;
    reg node462;
    reg node463;
    reg node464_r;
    reg node464_l;
    reg node465_r;
    reg node465_l;
    reg node466_r;
    reg node466_l;
    reg node467;
    reg node468;
    reg node469_r;
    reg node469_l;
    reg node470;
    reg node471;
    reg node472_r;
    reg node472_l;
    reg node473_r;
    reg node473_l;
    reg node474;
    reg node475;
    reg node476_r;
    reg node476_l;
    reg node477;
    reg node478;
    reg node479_r;
    reg node479_l;
    reg node480_r;
    reg node480_l;
    reg node481_r;
    reg node481_l;
    reg node482_r;
    reg node482_l;
    reg node483_r;
    reg node483_l;
    reg node484;
    reg node485;
    reg node486_r;
    reg node486_l;
    reg node487;
    reg node488;
    reg node489_r;
    reg node489_l;
    reg node490_r;
    reg node490_l;
    reg node491;
    reg node492;
    reg node493_r;
    reg node493_l;
    reg node494;
    reg node495;
    reg node496_r;
    reg node496_l;
    reg node497_r;
    reg node497_l;
    reg node498_r;
    reg node498_l;
    reg node499;
    reg node500;
    reg node501_r;
    reg node501_l;
    reg node502;
    reg node503;
    reg node504_r;
    reg node504_l;
    reg node505_r;
    reg node505_l;
    reg node506;
    reg node507;
    reg node508_r;
    reg node508_l;
    reg node509;
    reg node510;
    reg node511_r;
    reg node511_l;
    reg node512_r;
    reg node512_l;
    reg node513_r;
    reg node513_l;
    reg node514_r;
    reg node514_l;
    reg node515;
    reg node516;
    reg node517_r;
    reg node517_l;
    reg node518;
    reg node519;
    reg node520_r;
    reg node520_l;
    reg node521_r;
    reg node521_l;
    reg node522;
    reg node523;
    reg node524_r;
    reg node524_l;
    reg node525;
    reg node526;
    reg node527_r;
    reg node527_l;
    reg node528_r;
    reg node528_l;
    reg node529_r;
    reg node529_l;
    reg node530;
    reg node531;
    reg node532;
    reg node533_r;
    reg node533_l;
    reg node534_r;
    reg node534_l;
    reg node535;
    reg node536;
    reg node537_r;
    reg node537_l;
    reg node538;
    reg node539;
    reg node540_r;
    reg node540_l;
    reg node541_r;
    reg node541_l;
    reg node542_r;
    reg node542_l;
    reg node543_r;
    reg node543_l;
    reg node544_r;
    reg node544_l;
    reg node545_r;
    reg node545_l;
    reg node546;
    reg node547;
    reg node548_r;
    reg node548_l;
    reg node549;
    reg node550;
    reg node551_r;
    reg node551_l;
    reg node552_r;
    reg node552_l;
    reg node553;
    reg node554;
    reg node555_r;
    reg node555_l;
    reg node556;
    reg node557;
    reg node558_r;
    reg node558_l;
    reg node559_r;
    reg node559_l;
    reg node560_r;
    reg node560_l;
    reg node561;
    reg node562;
    reg node563_r;
    reg node563_l;
    reg node564;
    reg node565;
    reg node566_r;
    reg node566_l;
    reg node567_r;
    reg node567_l;
    reg node568;
    reg node569;
    reg node570_r;
    reg node570_l;
    reg node571;
    reg node572;
    reg node573_r;
    reg node573_l;
    reg node574_r;
    reg node574_l;
    reg node575_r;
    reg node575_l;
    reg node576_r;
    reg node576_l;
    reg node577;
    reg node578;
    reg node579_r;
    reg node579_l;
    reg node580;
    reg node581;
    reg node582_r;
    reg node582_l;
    reg node583_r;
    reg node583_l;
    reg node584;
    reg node585;
    reg node586_r;
    reg node586_l;
    reg node587;
    reg node588;
    reg node589;
    reg node590_r;
    reg node590_l;
    reg node591_r;
    reg node591_l;
    reg node592_r;
    reg node592_l;
    reg node593;
    reg node594_r;
    reg node594_l;
    reg node595;
    reg node596;
    reg node597_r;
    reg node597_l;
    reg node598;
    reg node599;
    reg node600_r;
    reg node600_l;
    reg node601_r;
    reg node601_l;
    reg node602_r;
    reg node602_l;
    reg node603;
    reg node604;
    reg node605;
    reg node606_r;
    reg node606_l;
    reg node607;
    reg node608_r;
    reg node608_l;
    reg node609;
    reg node610;
    reg node611_r;
    reg node611_l;
    reg node612_r;
    reg node612_l;
    reg node613_r;
    reg node613_l;
    reg node614_r;
    reg node614_l;
    reg node615_r;
    reg node615_l;
    reg node616_r;
    reg node616_l;
    reg node617_r;
    reg node617_l;
    reg node618;
    reg node619;
    reg node620_r;
    reg node620_l;
    reg node621;
    reg node622;
    reg node623_r;
    reg node623_l;
    reg node624_r;
    reg node624_l;
    reg node625;
    reg node626;
    reg node627_r;
    reg node627_l;
    reg node628;
    reg node629;
    reg node630_r;
    reg node630_l;
    reg node631_r;
    reg node631_l;
    reg node632_r;
    reg node632_l;
    reg node633;
    reg node634;
    reg node635_r;
    reg node635_l;
    reg node636;
    reg node637;
    reg node638_r;
    reg node638_l;
    reg node639_r;
    reg node639_l;
    reg node640;
    reg node641;
    reg node642;
    reg node643_r;
    reg node643_l;
    reg node644_r;
    reg node644_l;
    reg node645_r;
    reg node645_l;
    reg node646_r;
    reg node646_l;
    reg node647;
    reg node648;
    reg node649;
    reg node650_r;
    reg node650_l;
    reg node651;
    reg node652_r;
    reg node652_l;
    reg node653;
    reg node654;
    reg node655_r;
    reg node655_l;
    reg node656;
    reg node657;
    reg node658_r;
    reg node658_l;
    reg node659_r;
    reg node659_l;
    reg node660_r;
    reg node660_l;
    reg node661_r;
    reg node661_l;
    reg node662_r;
    reg node662_l;
    reg node663;
    reg node664;
    reg node665_r;
    reg node665_l;
    reg node666;
    reg node667;
    reg node668_r;
    reg node668_l;
    reg node669_r;
    reg node669_l;
    reg node670;
    reg node671;
    reg node672_r;
    reg node672_l;
    reg node673;
    reg node674;
    reg node675_r;
    reg node675_l;
    reg node676_r;
    reg node676_l;
    reg node677_r;
    reg node677_l;
    reg node678;
    reg node679;
    reg node680_r;
    reg node680_l;
    reg node681;
    reg node682;
    reg node683_r;
    reg node683_l;
    reg node684_r;
    reg node684_l;
    reg node685;
    reg node686;
    reg node687_r;
    reg node687_l;
    reg node688;
    reg node689;
    reg node690_r;
    reg node690_l;
    reg node691_r;
    reg node691_l;
    reg node692_r;
    reg node692_l;
    reg node693_r;
    reg node693_l;
    reg node694;
    reg node695;
    reg node696_r;
    reg node696_l;
    reg node697;
    reg node698;
    reg node699_r;
    reg node699_l;
    reg node700;
    reg node701;
    reg node702_r;
    reg node702_l;
    reg node703_r;
    reg node703_l;
    reg node704_r;
    reg node704_l;
    reg node705;
    reg node706;
    reg node707_r;
    reg node707_l;
    reg node708;
    reg node709;
    reg node710_r;
    reg node710_l;
    reg node711_r;
    reg node711_l;
    reg node712;
    reg node713;
    reg node714;
    reg node715_r;
    reg node715_l;
    reg node716_r;
    reg node716_l;
    reg node717_r;
    reg node717_l;
    reg node718_r;
    reg node718_l;
    reg node719_r;
    reg node719_l;
    reg node720_r;
    reg node720_l;
    reg node721;
    reg node722;
    reg node723_r;
    reg node723_l;
    reg node724;
    reg node725;
    reg node726_r;
    reg node726_l;
    reg node727_r;
    reg node727_l;
    reg node728;
    reg node729;
    reg node730_r;
    reg node730_l;
    reg node731;
    reg node732;
    reg node733_r;
    reg node733_l;
    reg node734_r;
    reg node734_l;
    reg node735_r;
    reg node735_l;
    reg node736;
    reg node737;
    reg node738_r;
    reg node738_l;
    reg node739;
    reg node740;
    reg node741_r;
    reg node741_l;
    reg node742_r;
    reg node742_l;
    reg node743;
    reg node744;
    reg node745_r;
    reg node745_l;
    reg node746;
    reg node747;
    reg node748_r;
    reg node748_l;
    reg node749_r;
    reg node749_l;
    reg node750_r;
    reg node750_l;
    reg node751_r;
    reg node751_l;
    reg node752;
    reg node753;
    reg node754_r;
    reg node754_l;
    reg node755;
    reg node756;
    reg node757_r;
    reg node757_l;
    reg node758_r;
    reg node758_l;
    reg node759;
    reg node760;
    reg node761_r;
    reg node761_l;
    reg node762;
    reg node763;
    reg node764_r;
    reg node764_l;
    reg node765_r;
    reg node765_l;
    reg node766_r;
    reg node766_l;
    reg node767;
    reg node768;
    reg node769;
    reg node770_r;
    reg node770_l;
    reg node771_r;
    reg node771_l;
    reg node772;
    reg node773;
    reg node774_r;
    reg node774_l;
    reg node775;
    reg node776;
    reg node777_r;
    reg node777_l;
    reg node778_r;
    reg node778_l;
    reg node779_r;
    reg node779_l;
    reg node780_r;
    reg node780_l;
    reg node781_r;
    reg node781_l;
    reg node782;
    reg node783;
    reg node784_r;
    reg node784_l;
    reg node785;
    reg node786;
    reg node787_r;
    reg node787_l;
    reg node788_r;
    reg node788_l;
    reg node789;
    reg node790;
    reg node791_r;
    reg node791_l;
    reg node792;
    reg node793;
    reg node794_r;
    reg node794_l;
    reg node795_r;
    reg node795_l;
    reg node796_r;
    reg node796_l;
    reg node797;
    reg node798;
    reg node799_r;
    reg node799_l;
    reg node800;
    reg node801;
    reg node802;
    reg node803_r;
    reg node803_l;
    reg node804_r;
    reg node804_l;
    reg node805_r;
    reg node805_l;
    reg node806;
    reg node807;
    reg node808_r;
    reg node808_l;
    reg node809;
    reg node810;
    reg node811_r;
    reg node811_l;
    reg node812;
    reg node813_r;
    reg node813_l;
    reg node814;
    reg node815;
    reg node816_r;
    reg node816_l;
    reg node817_r;
    reg node817_l;
    reg node818_r;
    reg node818_l;
    reg node819_r;
    reg node819_l;
    reg node820_r;
    reg node820_l;
    reg node821_r;
    reg node821_l;
    reg node822_r;
    reg node822_l;
    reg node823_r;
    reg node823_l;
    reg node824_r;
    reg node824_l;
    reg node825;
    reg node826;
    reg node827_r;
    reg node827_l;
    reg node828;
    reg node829;
    reg node830_r;
    reg node830_l;
    reg node831_r;
    reg node831_l;
    reg node832;
    reg node833;
    reg node834_r;
    reg node834_l;
    reg node835;
    reg node836;
    reg node837_r;
    reg node837_l;
    reg node838_r;
    reg node838_l;
    reg node839_r;
    reg node839_l;
    reg node840;
    reg node841;
    reg node842_r;
    reg node842_l;
    reg node843;
    reg node844;
    reg node845_r;
    reg node845_l;
    reg node846_r;
    reg node846_l;
    reg node847;
    reg node848;
    reg node849_r;
    reg node849_l;
    reg node850;
    reg node851;
    reg node852_r;
    reg node852_l;
    reg node853_r;
    reg node853_l;
    reg node854_r;
    reg node854_l;
    reg node855_r;
    reg node855_l;
    reg node856;
    reg node857;
    reg node858_r;
    reg node858_l;
    reg node859;
    reg node860;
    reg node861_r;
    reg node861_l;
    reg node862_r;
    reg node862_l;
    reg node863;
    reg node864;
    reg node865_r;
    reg node865_l;
    reg node866;
    reg node867;
    reg node868_r;
    reg node868_l;
    reg node869_r;
    reg node869_l;
    reg node870_r;
    reg node870_l;
    reg node871;
    reg node872;
    reg node873_r;
    reg node873_l;
    reg node874;
    reg node875;
    reg node876_r;
    reg node876_l;
    reg node877_r;
    reg node877_l;
    reg node878;
    reg node879;
    reg node880_r;
    reg node880_l;
    reg node881;
    reg node882;
    reg node883_r;
    reg node883_l;
    reg node884_r;
    reg node884_l;
    reg node885_r;
    reg node885_l;
    reg node886_r;
    reg node886_l;
    reg node887;
    reg node888;
    reg node889_r;
    reg node889_l;
    reg node890_r;
    reg node890_l;
    reg node891;
    reg node892;
    reg node893_r;
    reg node893_l;
    reg node894;
    reg node895;
    reg node896;
    reg node897_r;
    reg node897_l;
    reg node898_r;
    reg node898_l;
    reg node899_r;
    reg node899_l;
    reg node900_r;
    reg node900_l;
    reg node901;
    reg node902;
    reg node903_r;
    reg node903_l;
    reg node904;
    reg node905;
    reg node906_r;
    reg node906_l;
    reg node907_r;
    reg node907_l;
    reg node908;
    reg node909;
    reg node910_r;
    reg node910_l;
    reg node911;
    reg node912;
    reg node913_r;
    reg node913_l;
    reg node914_r;
    reg node914_l;
    reg node915_r;
    reg node915_l;
    reg node916;
    reg node917;
    reg node918_r;
    reg node918_l;
    reg node919;
    reg node920;
    reg node921_r;
    reg node921_l;
    reg node922_r;
    reg node922_l;
    reg node923;
    reg node924;
    reg node925_r;
    reg node925_l;
    reg node926;
    reg node927;
    reg node928_r;
    reg node928_l;
    reg node929_r;
    reg node929_l;
    reg node930_r;
    reg node930_l;
    reg node931_r;
    reg node931_l;
    reg node932_r;
    reg node932_l;
    reg node933_r;
    reg node933_l;
    reg node934;
    reg node935;
    reg node936_r;
    reg node936_l;
    reg node937;
    reg node938;
    reg node939_r;
    reg node939_l;
    reg node940_r;
    reg node940_l;
    reg node941;
    reg node942;
    reg node943_r;
    reg node943_l;
    reg node944;
    reg node945;
    reg node946_r;
    reg node946_l;
    reg node947_r;
    reg node947_l;
    reg node948_r;
    reg node948_l;
    reg node949;
    reg node950;
    reg node951_r;
    reg node951_l;
    reg node952;
    reg node953;
    reg node954_r;
    reg node954_l;
    reg node955_r;
    reg node955_l;
    reg node956;
    reg node957;
    reg node958_r;
    reg node958_l;
    reg node959;
    reg node960;
    reg node961_r;
    reg node961_l;
    reg node962_r;
    reg node962_l;
    reg node963_r;
    reg node963_l;
    reg node964_r;
    reg node964_l;
    reg node965;
    reg node966;
    reg node967;
    reg node968_r;
    reg node968_l;
    reg node969_r;
    reg node969_l;
    reg node970;
    reg node971;
    reg node972;
    reg node973_r;
    reg node973_l;
    reg node974_r;
    reg node974_l;
    reg node975_r;
    reg node975_l;
    reg node976;
    reg node977;
    reg node978;
    reg node979_r;
    reg node979_l;
    reg node980_r;
    reg node980_l;
    reg node981;
    reg node982;
    reg node983_r;
    reg node983_l;
    reg node984;
    reg node985;
    reg node986_r;
    reg node986_l;
    reg node987_r;
    reg node987_l;
    reg node988_r;
    reg node988_l;
    reg node989_r;
    reg node989_l;
    reg node990_r;
    reg node990_l;
    reg node991;
    reg node992;
    reg node993_r;
    reg node993_l;
    reg node994;
    reg node995;
    reg node996_r;
    reg node996_l;
    reg node997_r;
    reg node997_l;
    reg node998;
    reg node999;
    reg node1000_r;
    reg node1000_l;
    reg node1001;
    reg node1002;
    reg node1003_r;
    reg node1003_l;
    reg node1004_r;
    reg node1004_l;
    reg node1005_r;
    reg node1005_l;
    reg node1006;
    reg node1007;
    reg node1008_r;
    reg node1008_l;
    reg node1009;
    reg node1010;
    reg node1011_r;
    reg node1011_l;
    reg node1012_r;
    reg node1012_l;
    reg node1013;
    reg node1014;
    reg node1015_r;
    reg node1015_l;
    reg node1016;
    reg node1017;
    reg node1018_r;
    reg node1018_l;
    reg node1019_r;
    reg node1019_l;
    reg node1020_r;
    reg node1020_l;
    reg node1021_r;
    reg node1021_l;
    reg node1022;
    reg node1023;
    reg node1024_r;
    reg node1024_l;
    reg node1025;
    reg node1026;
    reg node1027_r;
    reg node1027_l;
    reg node1028_r;
    reg node1028_l;
    reg node1029;
    reg node1030;
    reg node1031_r;
    reg node1031_l;
    reg node1032;
    reg node1033;
    reg node1034_r;
    reg node1034_l;
    reg node1035_r;
    reg node1035_l;
    reg node1036_r;
    reg node1036_l;
    reg node1037;
    reg node1038;
    reg node1039_r;
    reg node1039_l;
    reg node1040;
    reg node1041;
    reg node1042_r;
    reg node1042_l;
    reg node1043_r;
    reg node1043_l;
    reg node1044;
    reg node1045;
    reg node1046_r;
    reg node1046_l;
    reg node1047;
    reg node1048;
    reg node1049_r;
    reg node1049_l;
    reg node1050_r;
    reg node1050_l;
    reg node1051_r;
    reg node1051_l;
    reg node1052_r;
    reg node1052_l;
    reg node1053_r;
    reg node1053_l;
    reg node1054_r;
    reg node1054_l;
    reg node1055_r;
    reg node1055_l;
    reg node1056;
    reg node1057;
    reg node1058_r;
    reg node1058_l;
    reg node1059;
    reg node1060;
    reg node1061_r;
    reg node1061_l;
    reg node1062_r;
    reg node1062_l;
    reg node1063;
    reg node1064;
    reg node1065;
    reg node1066_r;
    reg node1066_l;
    reg node1067_r;
    reg node1067_l;
    reg node1068_r;
    reg node1068_l;
    reg node1069;
    reg node1070;
    reg node1071;
    reg node1072_r;
    reg node1072_l;
    reg node1073_r;
    reg node1073_l;
    reg node1074;
    reg node1075;
    reg node1076_r;
    reg node1076_l;
    reg node1077;
    reg node1078;
    reg node1079_r;
    reg node1079_l;
    reg node1080_r;
    reg node1080_l;
    reg node1081_r;
    reg node1081_l;
    reg node1082_r;
    reg node1082_l;
    reg node1083;
    reg node1084;
    reg node1085_r;
    reg node1085_l;
    reg node1086;
    reg node1087;
    reg node1088_r;
    reg node1088_l;
    reg node1089;
    reg node1090_r;
    reg node1090_l;
    reg node1091;
    reg node1092;
    reg node1093_r;
    reg node1093_l;
    reg node1094_r;
    reg node1094_l;
    reg node1095_r;
    reg node1095_l;
    reg node1096;
    reg node1097;
    reg node1098_r;
    reg node1098_l;
    reg node1099;
    reg node1100;
    reg node1101_r;
    reg node1101_l;
    reg node1102_r;
    reg node1102_l;
    reg node1103;
    reg node1104;
    reg node1105_r;
    reg node1105_l;
    reg node1106;
    reg node1107;
    reg node1108_r;
    reg node1108_l;
    reg node1109_r;
    reg node1109_l;
    reg node1110_r;
    reg node1110_l;
    reg node1111_r;
    reg node1111_l;
    reg node1112_r;
    reg node1112_l;
    reg node1113;
    reg node1114;
    reg node1115_r;
    reg node1115_l;
    reg node1116;
    reg node1117;
    reg node1118_r;
    reg node1118_l;
    reg node1119_r;
    reg node1119_l;
    reg node1120;
    reg node1121;
    reg node1122_r;
    reg node1122_l;
    reg node1123;
    reg node1124;
    reg node1125_r;
    reg node1125_l;
    reg node1126_r;
    reg node1126_l;
    reg node1127_r;
    reg node1127_l;
    reg node1128;
    reg node1129;
    reg node1130_r;
    reg node1130_l;
    reg node1131;
    reg node1132;
    reg node1133_r;
    reg node1133_l;
    reg node1134_r;
    reg node1134_l;
    reg node1135;
    reg node1136;
    reg node1137_r;
    reg node1137_l;
    reg node1138;
    reg node1139;
    reg node1140_r;
    reg node1140_l;
    reg node1141_r;
    reg node1141_l;
    reg node1142_r;
    reg node1142_l;
    reg node1143_r;
    reg node1143_l;
    reg node1144;
    reg node1145;
    reg node1146_r;
    reg node1146_l;
    reg node1147;
    reg node1148;
    reg node1149_r;
    reg node1149_l;
    reg node1150_r;
    reg node1150_l;
    reg node1151;
    reg node1152;
    reg node1153_r;
    reg node1153_l;
    reg node1154;
    reg node1155;
    reg node1156_r;
    reg node1156_l;
    reg node1157_r;
    reg node1157_l;
    reg node1158_r;
    reg node1158_l;
    reg node1159;
    reg node1160;
    reg node1161_r;
    reg node1161_l;
    reg node1162;
    reg node1163;
    reg node1164_r;
    reg node1164_l;
    reg node1165_r;
    reg node1165_l;
    reg node1166;
    reg node1167;
    reg node1168_r;
    reg node1168_l;
    reg node1169;
    reg node1170;
    reg node1171_r;
    reg node1171_l;
    reg node1172_r;
    reg node1172_l;
    reg node1173_r;
    reg node1173_l;
    reg node1174_r;
    reg node1174_l;
    reg node1175_r;
    reg node1175_l;
    reg node1176_r;
    reg node1176_l;
    reg node1177;
    reg node1178;
    reg node1179_r;
    reg node1179_l;
    reg node1180;
    reg node1181;
    reg node1182_r;
    reg node1182_l;
    reg node1183_r;
    reg node1183_l;
    reg node1184;
    reg node1185;
    reg node1186_r;
    reg node1186_l;
    reg node1187;
    reg node1188;
    reg node1189_r;
    reg node1189_l;
    reg node1190_r;
    reg node1190_l;
    reg node1191_r;
    reg node1191_l;
    reg node1192;
    reg node1193;
    reg node1194_r;
    reg node1194_l;
    reg node1195;
    reg node1196;
    reg node1197_r;
    reg node1197_l;
    reg node1198;
    reg node1199;
    reg node1200_r;
    reg node1200_l;
    reg node1201_r;
    reg node1201_l;
    reg node1202;
    reg node1203_r;
    reg node1203_l;
    reg node1204;
    reg node1205;
    reg node1206_r;
    reg node1206_l;
    reg node1207;
    reg node1208_r;
    reg node1208_l;
    reg node1209_r;
    reg node1209_l;
    reg node1210;
    reg node1211;
    reg node1212;
    reg node1213_r;
    reg node1213_l;
    reg node1214_r;
    reg node1214_l;
    reg node1215_r;
    reg node1215_l;
    reg node1216_r;
    reg node1216_l;
    reg node1217_r;
    reg node1217_l;
    reg node1218;
    reg node1219;
    reg node1220_r;
    reg node1220_l;
    reg node1221;
    reg node1222;
    reg node1223_r;
    reg node1223_l;
    reg node1224_r;
    reg node1224_l;
    reg node1225;
    reg node1226;
    reg node1227_r;
    reg node1227_l;
    reg node1228;
    reg node1229;
    reg node1230_r;
    reg node1230_l;
    reg node1231_r;
    reg node1231_l;
    reg node1232_r;
    reg node1232_l;
    reg node1233;
    reg node1234;
    reg node1235_r;
    reg node1235_l;
    reg node1236;
    reg node1237;
    reg node1238_r;
    reg node1238_l;
    reg node1239_r;
    reg node1239_l;
    reg node1240;
    reg node1241;
    reg node1242_r;
    reg node1242_l;
    reg node1243;
    reg node1244;
    reg node1245_r;
    reg node1245_l;
    reg node1246_r;
    reg node1246_l;
    reg node1247_r;
    reg node1247_l;
    reg node1248_r;
    reg node1248_l;
    reg node1249;
    reg node1250;
    reg node1251_r;
    reg node1251_l;
    reg node1252;
    reg node1253;
    reg node1254_r;
    reg node1254_l;
    reg node1255_r;
    reg node1255_l;
    reg node1256;
    reg node1257;
    reg node1258;
    reg node1259_r;
    reg node1259_l;
    reg node1260_r;
    reg node1260_l;
    reg node1261_r;
    reg node1261_l;
    reg node1262;
    reg node1263;
    reg node1264_r;
    reg node1264_l;
    reg node1265;
    reg node1266;
    reg node1267_r;
    reg node1267_l;
    reg node1268_r;
    reg node1268_l;
    reg node1269;
    reg node1270;
    reg node1271_r;
    reg node1271_l;
    reg node1272;
    reg node1273;
    reg node1274_r;
    reg node1274_l;
    reg node1275_r;
    reg node1275_l;
    reg node1276_r;
    reg node1276_l;
    reg node1277_r;
    reg node1277_l;
    reg node1278_r;
    reg node1278_l;
    reg node1279_r;
    reg node1279_l;
    reg node1280_r;
    reg node1280_l;
    reg node1281_r;
    reg node1281_l;
    reg node1282;
    reg node1283;
    reg node1284_r;
    reg node1284_l;
    reg node1285;
    reg node1286;
    reg node1287_r;
    reg node1287_l;
    reg node1288_r;
    reg node1288_l;
    reg node1289;
    reg node1290;
    reg node1291_r;
    reg node1291_l;
    reg node1292;
    reg node1293;
    reg node1294_r;
    reg node1294_l;
    reg node1295_r;
    reg node1295_l;
    reg node1296_r;
    reg node1296_l;
    reg node1297;
    reg node1298;
    reg node1299_r;
    reg node1299_l;
    reg node1300;
    reg node1301;
    reg node1302_r;
    reg node1302_l;
    reg node1303_r;
    reg node1303_l;
    reg node1304;
    reg node1305;
    reg node1306_r;
    reg node1306_l;
    reg node1307;
    reg node1308;
    reg node1309_r;
    reg node1309_l;
    reg node1310_r;
    reg node1310_l;
    reg node1311_r;
    reg node1311_l;
    reg node1312_r;
    reg node1312_l;
    reg node1313;
    reg node1314;
    reg node1315_r;
    reg node1315_l;
    reg node1316;
    reg node1317;
    reg node1318_r;
    reg node1318_l;
    reg node1319_r;
    reg node1319_l;
    reg node1320;
    reg node1321;
    reg node1322_r;
    reg node1322_l;
    reg node1323;
    reg node1324;
    reg node1325_r;
    reg node1325_l;
    reg node1326_r;
    reg node1326_l;
    reg node1327_r;
    reg node1327_l;
    reg node1328;
    reg node1329;
    reg node1330_r;
    reg node1330_l;
    reg node1331;
    reg node1332;
    reg node1333_r;
    reg node1333_l;
    reg node1334_r;
    reg node1334_l;
    reg node1335;
    reg node1336;
    reg node1337_r;
    reg node1337_l;
    reg node1338;
    reg node1339;
    reg node1340_r;
    reg node1340_l;
    reg node1341_r;
    reg node1341_l;
    reg node1342_r;
    reg node1342_l;
    reg node1343_r;
    reg node1343_l;
    reg node1344_r;
    reg node1344_l;
    reg node1345;
    reg node1346;
    reg node1347;
    reg node1348_r;
    reg node1348_l;
    reg node1349_r;
    reg node1349_l;
    reg node1350;
    reg node1351;
    reg node1352_r;
    reg node1352_l;
    reg node1353;
    reg node1354;
    reg node1355_r;
    reg node1355_l;
    reg node1356_r;
    reg node1356_l;
    reg node1357;
    reg node1358;
    reg node1359;
    reg node1360_r;
    reg node1360_l;
    reg node1361_r;
    reg node1361_l;
    reg node1362_r;
    reg node1362_l;
    reg node1363_r;
    reg node1363_l;
    reg node1364;
    reg node1365;
    reg node1366_r;
    reg node1366_l;
    reg node1367;
    reg node1368;
    reg node1369_r;
    reg node1369_l;
    reg node1370_r;
    reg node1370_l;
    reg node1371;
    reg node1372;
    reg node1373;
    reg node1374_r;
    reg node1374_l;
    reg node1375_r;
    reg node1375_l;
    reg node1376;
    reg node1377_r;
    reg node1377_l;
    reg node1378;
    reg node1379;
    reg node1380_r;
    reg node1380_l;
    reg node1381_r;
    reg node1381_l;
    reg node1382;
    reg node1383;
    reg node1384_r;
    reg node1384_l;
    reg node1385;
    reg node1386;
    reg node1387_r;
    reg node1387_l;
    reg node1388_r;
    reg node1388_l;
    reg node1389_r;
    reg node1389_l;
    reg node1390_r;
    reg node1390_l;
    reg node1391_r;
    reg node1391_l;
    reg node1392;
    reg node1393_r;
    reg node1393_l;
    reg node1394;
    reg node1395;
    reg node1396_r;
    reg node1396_l;
    reg node1397_r;
    reg node1397_l;
    reg node1398;
    reg node1399;
    reg node1400_r;
    reg node1400_l;
    reg node1401;
    reg node1402;
    reg node1403_r;
    reg node1403_l;
    reg node1404;
    reg node1405_r;
    reg node1405_l;
    reg node1406_r;
    reg node1406_l;
    reg node1407;
    reg node1408;
    reg node1409;
    reg node1410_r;
    reg node1410_l;
    reg node1411_r;
    reg node1411_l;
    reg node1412_r;
    reg node1412_l;
    reg node1413_r;
    reg node1413_l;
    reg node1414;
    reg node1415;
    reg node1416_r;
    reg node1416_l;
    reg node1417;
    reg node1418;
    reg node1419_r;
    reg node1419_l;
    reg node1420_r;
    reg node1420_l;
    reg node1421;
    reg node1422;
    reg node1423_r;
    reg node1423_l;
    reg node1424;
    reg node1425;
    reg node1426_r;
    reg node1426_l;
    reg node1427_r;
    reg node1427_l;
    reg node1428_r;
    reg node1428_l;
    reg node1429;
    reg node1430;
    reg node1431;
    reg node1432_r;
    reg node1432_l;
    reg node1433_r;
    reg node1433_l;
    reg node1434;
    reg node1435;
    reg node1436;
    reg node1437_r;
    reg node1437_l;
    reg node1438_r;
    reg node1438_l;
    reg node1439_r;
    reg node1439_l;
    reg node1440_r;
    reg node1440_l;
    reg node1441_r;
    reg node1441_l;
    reg node1442;
    reg node1443;
    reg node1444_r;
    reg node1444_l;
    reg node1445;
    reg node1446;
    reg node1447_r;
    reg node1447_l;
    reg node1448_r;
    reg node1448_l;
    reg node1449;
    reg node1450;
    reg node1451_r;
    reg node1451_l;
    reg node1452;
    reg node1453;
    reg node1454_r;
    reg node1454_l;
    reg node1455_r;
    reg node1455_l;
    reg node1456_r;
    reg node1456_l;
    reg node1457;
    reg node1458;
    reg node1459_r;
    reg node1459_l;
    reg node1460;
    reg node1461;
    reg node1462_r;
    reg node1462_l;
    reg node1463_r;
    reg node1463_l;
    reg node1464;
    reg node1465;
    reg node1466_r;
    reg node1466_l;
    reg node1467;
    reg node1468;
    reg node1469_r;
    reg node1469_l;
    reg node1470_r;
    reg node1470_l;
    reg node1471_r;
    reg node1471_l;
    reg node1472_r;
    reg node1472_l;
    reg node1473;
    reg node1474;
    reg node1475_r;
    reg node1475_l;
    reg node1476;
    reg node1477;
    reg node1478_r;
    reg node1478_l;
    reg node1479_r;
    reg node1479_l;
    reg node1480;
    reg node1481;
    reg node1482_r;
    reg node1482_l;
    reg node1483;
    reg node1484;
    reg node1485_r;
    reg node1485_l;
    reg node1486_r;
    reg node1486_l;
    reg node1487_r;
    reg node1487_l;
    reg node1488;
    reg node1489;
    reg node1490_r;
    reg node1490_l;
    reg node1491;
    reg node1492;
    reg node1493_r;
    reg node1493_l;
    reg node1494_r;
    reg node1494_l;
    reg node1495;
    reg node1496;
    reg node1497_r;
    reg node1497_l;
    reg node1498;
    reg node1499;
    reg node1500_r;
    reg node1500_l;
    reg node1501_r;
    reg node1501_l;
    reg node1502_r;
    reg node1502_l;
    reg node1503_r;
    reg node1503_l;
    reg node1504_r;
    reg node1504_l;
    reg node1505_r;
    reg node1505_l;
    reg node1506_r;
    reg node1506_l;
    reg node1507;
    reg node1508;
    reg node1509;
    reg node1510_r;
    reg node1510_l;
    reg node1511;
    reg node1512;
    reg node1513_r;
    reg node1513_l;
    reg node1514_r;
    reg node1514_l;
    reg node1515_r;
    reg node1515_l;
    reg node1516;
    reg node1517;
    reg node1518;
    reg node1519_r;
    reg node1519_l;
    reg node1520_r;
    reg node1520_l;
    reg node1521;
    reg node1522;
    reg node1523_r;
    reg node1523_l;
    reg node1524;
    reg node1525;
    reg node1526_r;
    reg node1526_l;
    reg node1527_r;
    reg node1527_l;
    reg node1528_r;
    reg node1528_l;
    reg node1529_r;
    reg node1529_l;
    reg node1530;
    reg node1531;
    reg node1532_r;
    reg node1532_l;
    reg node1533;
    reg node1534;
    reg node1535_r;
    reg node1535_l;
    reg node1536_r;
    reg node1536_l;
    reg node1537;
    reg node1538;
    reg node1539;
    reg node1540_r;
    reg node1540_l;
    reg node1541_r;
    reg node1541_l;
    reg node1542_r;
    reg node1542_l;
    reg node1543;
    reg node1544;
    reg node1545;
    reg node1546_r;
    reg node1546_l;
    reg node1547_r;
    reg node1547_l;
    reg node1548;
    reg node1549;
    reg node1550_r;
    reg node1550_l;
    reg node1551;
    reg node1552;
    reg node1553_r;
    reg node1553_l;
    reg node1554_r;
    reg node1554_l;
    reg node1555;
    reg node1556_r;
    reg node1556_l;
    reg node1557_r;
    reg node1557_l;
    reg node1558;
    reg node1559_r;
    reg node1559_l;
    reg node1560;
    reg node1561;
    reg node1562;
    reg node1563_r;
    reg node1563_l;
    reg node1564;
    reg node1565;
    reg node1566_r;
    reg node1566_l;
    reg node1567_r;
    reg node1567_l;
    reg node1568_r;
    reg node1568_l;
    reg node1569_r;
    reg node1569_l;
    reg node1570;
    reg node1571;
    reg node1572_r;
    reg node1572_l;
    reg node1573;
    reg node1574_r;
    reg node1574_l;
    reg node1575;
    reg node1576_r;
    reg node1576_l;
    reg node1577;
    reg node1578;
    reg node1579_r;
    reg node1579_l;
    reg node1580_r;
    reg node1580_l;
    reg node1581;
    reg node1582;
    reg node1583_r;
    reg node1583_l;
    reg node1584_r;
    reg node1584_l;
    reg node1585_r;
    reg node1585_l;
    reg node1586;
    reg node1587;
    reg node1588;
    reg node1589_r;
    reg node1589_l;
    reg node1590;
    reg node1591;
    reg node1592_r;
    reg node1592_l;
    reg node1593_r;
    reg node1593_l;
    reg node1594_r;
    reg node1594_l;
    reg node1595_r;
    reg node1595_l;
    reg node1596;
    reg node1597_r;
    reg node1597_l;
    reg node1598;
    reg node1599;
    reg node1600_r;
    reg node1600_l;
    reg node1601;
    reg node1602;
    reg node1603_r;
    reg node1603_l;
    reg node1604_r;
    reg node1604_l;
    reg node1605_r;
    reg node1605_l;
    reg node1606;
    reg node1607;
    reg node1608_r;
    reg node1608_l;
    reg node1609;
    reg node1610;
    reg node1611_r;
    reg node1611_l;
    reg node1612;
    reg node1613_r;
    reg node1613_l;
    reg node1614;
    reg node1615;
    reg node1616_r;
    reg node1616_l;
    reg node1617_r;
    reg node1617_l;
    reg node1618_r;
    reg node1618_l;
    reg node1619;
    reg node1620;
    reg node1621;
    reg node1622_r;
    reg node1622_l;
    reg node1623_r;
    reg node1623_l;
    reg node1624;
    reg node1625_r;
    reg node1625_l;
    reg node1626;
    reg node1627;
    reg node1628_r;
    reg node1628_l;
    reg node1629_r;
    reg node1629_l;
    reg node1630;
    reg node1631;
    reg node1632;
    reg result0;
    reg result1;
    reg result2;
    reg result3;
    reg result4;
    reg result5;
    reg result6;
    reg result7;
    reg result8;
    reg result9;

    begin
      node0_r = pixel[409];
      node0_l = ~pixel[409];
      node1_r = node0_l & pixel[378];
      node1_l = node0_l & ~pixel[378];
      node2_r = node1_l & pixel[462];
      node2_l = node1_l & ~pixel[462];
      node3_r = node2_l & pixel[372];
      node3_l = node2_l & ~pixel[372];
      node4_r = node3_l & pixel[185];
      node4_l = node3_l & ~pixel[185];
      node5_r = node4_l & pixel[598];
      node5_l = node4_l & ~pixel[598];
      node6_r = node5_l & pixel[431];
      node6_l = node5_l & ~pixel[431];
      node7_r = node6_l & pixel[152];
      node7_l = node6_l & ~pixel[152];
      node8_r = node7_l & pixel[416];
      node8_l = node7_l & ~pixel[416];
      node9_r = node8_l & pixel[515];
      node9_l = node8_l & ~pixel[515];
      node10 = node9_l;
      node11 = node9_r;
      node12_r = node8_r & pixel[464];
      node12_l = node8_r & ~pixel[464];
      node13 = node12_l;
      node14 = node12_r;
      node15_r = node7_r & pixel[634];
      node15_l = node7_r & ~pixel[634];
      node16_r = node15_l & pixel[398];
      node16_l = node15_l & ~pixel[398];
      node17 = node16_l;
      node18 = node16_r;
      node19_r = node15_r & pixel[269];
      node19_l = node15_r & ~pixel[269];
      node20 = node19_l;
      node21 = node19_r;
      node22_r = node6_r & pixel[268];
      node22_l = node6_r & ~pixel[268];
      node23_r = node22_l & pixel[99];
      node23_l = node22_l & ~pixel[99];
      node24_r = node23_l & pixel[301];
      node24_l = node23_l & ~pixel[301];
      node25 = node24_l;
      node26 = node24_r;
      node27_r = node23_r & pixel[300];
      node27_l = node23_r & ~pixel[300];
      node28 = node27_l;
      node29 = node27_r;
      node30_r = node22_r & pixel[466];
      node30_l = node22_r & ~pixel[466];
      node31_r = node30_l & pixel[455];
      node31_l = node30_l & ~pixel[455];
      node32 = node31_l;
      node33 = node31_r;
      node34_r = node30_r & pixel[324];
      node34_l = node30_r & ~pixel[324];
      node35 = node34_l;
      node36 = node34_r;
      node37_r = node5_r & pixel[211];
      node37_l = node5_r & ~pixel[211];
      node38_r = node37_l & pixel[314];
      node38_l = node37_l & ~pixel[314];
      node39_r = node38_l & pixel[295];
      node39_l = node38_l & ~pixel[295];
      node40_r = node39_l & pixel[544];
      node40_l = node39_l & ~pixel[544];
      node41 = node40_l;
      node42 = node40_r;
      node43_r = node39_r & pixel[549];
      node43_l = node39_r & ~pixel[549];
      node44 = node43_l;
      node45 = node43_r;
      node46_r = node38_r & pixel[410];
      node46_l = node38_r & ~pixel[410];
      node47 = node46_l;
      node48_r = node46_r & pixel[354];
      node48_l = node46_r & ~pixel[354];
      node49 = node48_l;
      node50 = node48_r;
      node51_r = node37_r & pixel[454];
      node51_l = node37_r & ~pixel[454];
      node52_r = node51_l & pixel[345];
      node52_l = node51_l & ~pixel[345];
      node53_r = node52_l & pixel[263];
      node53_l = node52_l & ~pixel[263];
      node54 = node53_l;
      node55 = node53_r;
      node56_r = node52_r & pixel[353];
      node56_l = node52_r & ~pixel[353];
      node57 = node56_l;
      node58 = node56_r;
      node59_r = node51_r & pixel[212];
      node59_l = node51_r & ~pixel[212];
      node60 = node59_l;
      node61 = node59_r;
      node62_r = node4_r & pixel[401];
      node62_l = node4_r & ~pixel[401];
      node63_r = node62_l & pixel[481];
      node63_l = node62_l & ~pixel[481];
      node64_r = node63_l & pixel[430];
      node64_l = node63_l & ~pixel[430];
      node65_r = node64_l & pixel[324];
      node65_l = node64_l & ~pixel[324];
      node66_r = node65_l & pixel[546];
      node66_l = node65_l & ~pixel[546];
      node67 = node66_l;
      node68 = node66_r;
      node69_r = node65_r & pixel[263];
      node69_l = node65_r & ~pixel[263];
      node70 = node69_l;
      node71 = node69_r;
      node72_r = node64_r & pixel[411];
      node72_l = node64_r & ~pixel[411];
      node73_r = node72_l & pixel[656];
      node73_l = node72_l & ~pixel[656];
      node74 = node73_l;
      node75 = node73_r;
      node76_r = node72_r & pixel[490];
      node76_l = node72_r & ~pixel[490];
      node77 = node76_l;
      node78 = node76_r;
      node79_r = node63_r & pixel[323];
      node79_l = node63_r & ~pixel[323];
      node80_r = node79_l & pixel[489];
      node80_l = node79_l & ~pixel[489];
      node81_r = node80_l & pixel[638];
      node81_l = node80_l & ~pixel[638];
      node82 = node81_l;
      node83 = node81_r;
      node84_r = node80_r & pixel[608];
      node84_l = node80_r & ~pixel[608];
      node85 = node84_l;
      node86 = node84_r;
      node87_r = node79_r & pixel[315];
      node87_l = node79_r & ~pixel[315];
      node88_r = node87_l & pixel[122];
      node88_l = node87_l & ~pixel[122];
      node89 = node88_l;
      node90 = node88_r;
      node91 = node87_r;
      node92_r = node62_r & pixel[516];
      node92_l = node62_r & ~pixel[516];
      node93_r = node92_l & pixel[440];
      node93_l = node92_l & ~pixel[440];
      node94_r = node93_l & pixel[547];
      node94_l = node93_l & ~pixel[547];
      node95_r = node94_l & pixel[162];
      node95_l = node94_l & ~pixel[162];
      node96 = node95_l;
      node97 = node95_r;
      node98_r = node94_r & pixel[655];
      node98_l = node94_r & ~pixel[655];
      node99 = node98_l;
      node100 = node98_r;
      node101_r = node93_r & pixel[353];
      node101_l = node93_r & ~pixel[353];
      node102_r = node101_l & pixel[582];
      node102_l = node101_l & ~pixel[582];
      node103 = node102_l;
      node104 = node102_r;
      node105_r = node101_r & pixel[485];
      node105_l = node101_r & ~pixel[485];
      node106 = node105_l;
      node107 = node105_r;
      node108_r = node92_r & pixel[326];
      node108_l = node92_r & ~pixel[326];
      node109_r = node108_l & pixel[684];
      node109_l = node108_l & ~pixel[684];
      node110_r = node109_l & pixel[352];
      node110_l = node109_l & ~pixel[352];
      node111 = node110_l;
      node112 = node110_r;
      node113_r = node109_r & pixel[347];
      node113_l = node109_r & ~pixel[347];
      node114 = node113_l;
      node115 = node113_r;
      node116_r = node108_r & pixel[399];
      node116_l = node108_r & ~pixel[399];
      node117_r = node116_l & pixel[324];
      node117_l = node116_l & ~pixel[324];
      node118 = node117_l;
      node119 = node117_r;
      node120 = node116_r;
      node121_r = node3_r & pixel[483];
      node121_l = node3_r & ~pixel[483];
      node122_r = node121_l & pixel[480];
      node122_l = node121_l & ~pixel[480];
      node123_r = node122_l & pixel[512];
      node123_l = node122_l & ~pixel[512];
      node124_r = node123_l & pixel[383];
      node124_l = node123_l & ~pixel[383];
      node125_r = node124_l & pixel[454];
      node125_l = node124_l & ~pixel[454];
      node126_r = node125_l & pixel[553];
      node126_l = node125_l & ~pixel[553];
      node127 = node126_l;
      node128 = node126_r;
      node129_r = node125_r & pixel[510];
      node129_l = node125_r & ~pixel[510];
      node130 = node129_l;
      node131 = node129_r;
      node132_r = node124_r & pixel[513];
      node132_l = node124_r & ~pixel[513];
      node133_r = node132_l & pixel[322];
      node133_l = node132_l & ~pixel[322];
      node134 = node133_l;
      node135 = node133_r;
      node136_r = node132_r & pixel[376];
      node136_l = node132_r & ~pixel[376];
      node137 = node136_l;
      node138 = node136_r;
      node139_r = node123_r & pixel[328];
      node139_l = node123_r & ~pixel[328];
      node140_r = node139_l & pixel[487];
      node140_l = node139_l & ~pixel[487];
      node141_r = node140_l & pixel[221];
      node141_l = node140_l & ~pixel[221];
      node142 = node141_l;
      node143 = node141_r;
      node144_r = node140_r & pixel[573];
      node144_l = node140_r & ~pixel[573];
      node145 = node144_l;
      node146 = node144_r;
      node147_r = node139_r & pixel[272];
      node147_l = node139_r & ~pixel[272];
      node148_r = node147_l & pixel[295];
      node148_l = node147_l & ~pixel[295];
      node149 = node148_l;
      node150 = node148_r;
      node151_r = node147_r & pixel[648];
      node151_l = node147_r & ~pixel[648];
      node152 = node151_l;
      node153 = node151_r;
      node154_r = node122_r & pixel[509];
      node154_l = node122_r & ~pixel[509];
      node155_r = node154_l & pixel[565];
      node155_l = node154_l & ~pixel[565];
      node156 = node155_l;
      node157 = node155_r;
      node158_r = node154_r & pixel[459];
      node158_l = node154_r & ~pixel[459];
      node159_r = node158_l & pixel[375];
      node159_l = node158_l & ~pixel[375];
      node160_r = node159_l & pixel[689];
      node160_l = node159_l & ~pixel[689];
      node161 = node160_l;
      node162 = node160_r;
      node163_r = node159_r & pixel[358];
      node163_l = node159_r & ~pixel[358];
      node164 = node163_l;
      node165 = node163_r;
      node166_r = node158_r & pixel[492];
      node166_l = node158_r & ~pixel[492];
      node167 = node166_l;
      node168 = node166_r;
      node169_r = node121_r & pixel[716];
      node169_l = node121_r & ~pixel[716];
      node170_r = node169_l & pixel[597];
      node170_l = node169_l & ~pixel[597];
      node171_r = node170_l & pixel[715];
      node171_l = node170_l & ~pixel[715];
      node172_r = node171_l & pixel[492];
      node172_l = node171_l & ~pixel[492];
      node173_r = node172_l & pixel[690];
      node173_l = node172_l & ~pixel[690];
      node174 = node173_l;
      node175 = node173_r;
      node176_r = node172_r & pixel[636];
      node176_l = node172_r & ~pixel[636];
      node177 = node176_l;
      node178 = node176_r;
      node179 = node171_r;
      node180_r = node170_r & pixel[353];
      node180_l = node170_r & ~pixel[353];
      node181_r = node180_l & pixel[72];
      node181_l = node180_l & ~pixel[72];
      node182_r = node181_l & pixel[91];
      node182_l = node181_l & ~pixel[91];
      node183 = node182_l;
      node184 = node182_r;
      node185_r = node181_r & pixel[299];
      node185_l = node181_r & ~pixel[299];
      node186 = node185_l;
      node187 = node185_r;
      node188_r = node180_r & pixel[240];
      node188_l = node180_r & ~pixel[240];
      node189_r = node188_l & pixel[158];
      node189_l = node188_l & ~pixel[158];
      node190 = node189_l;
      node191 = node189_r;
      node192_r = node188_r & pixel[495];
      node192_l = node188_r & ~pixel[495];
      node193 = node192_l;
      node194 = node192_r;
      node195_r = node169_r & pixel[444];
      node195_l = node169_r & ~pixel[444];
      node196_r = node195_l & pixel[543];
      node196_l = node195_l & ~pixel[543];
      node197 = node196_l;
      node198_r = node196_r & pixel[383];
      node198_l = node196_r & ~pixel[383];
      node199 = node198_l;
      node200 = node198_r;
      node201 = node195_r;
      node202_r = node2_r & pixel[346];
      node202_l = node2_r & ~pixel[346];
      node203_r = node202_l & pixel[457];
      node203_l = node202_l & ~pixel[457];
      node204_r = node203_l & pixel[514];
      node204_l = node203_l & ~pixel[514];
      node205_r = node204_l & pixel[325];
      node205_l = node204_l & ~pixel[325];
      node206_r = node205_l & pixel[428];
      node206_l = node205_l & ~pixel[428];
      node207_r = node206_l & pixel[372];
      node207_l = node206_l & ~pixel[372];
      node208_r = node207_l & pixel[240];
      node208_l = node207_l & ~pixel[240];
      node209 = node208_l;
      node210 = node208_r;
      node211_r = node207_r & pixel[300];
      node211_l = node207_r & ~pixel[300];
      node212 = node211_l;
      node213 = node211_r;
      node214_r = node206_r & pixel[662];
      node214_l = node206_r & ~pixel[662];
      node215_r = node214_l & pixel[290];
      node215_l = node214_l & ~pixel[290];
      node216 = node215_l;
      node217 = node215_r;
      node218_r = node214_r & pixel[441];
      node218_l = node214_r & ~pixel[441];
      node219 = node218_l;
      node220 = node218_r;
      node221_r = node205_r & pixel[568];
      node221_l = node205_r & ~pixel[568];
      node222_r = node221_l & pixel[432];
      node222_l = node221_l & ~pixel[432];
      node223_r = node222_l & pixel[127];
      node223_l = node222_l & ~pixel[127];
      node224 = node223_l;
      node225 = node223_r;
      node226_r = node222_r & pixel[206];
      node226_l = node222_r & ~pixel[206];
      node227 = node226_l;
      node228 = node226_r;
      node229_r = node221_r & pixel[261];
      node229_l = node221_r & ~pixel[261];
      node230_r = node229_l & pixel[609];
      node230_l = node229_l & ~pixel[609];
      node231 = node230_l;
      node232 = node230_r;
      node233 = node229_r;
      node234_r = node204_r & pixel[241];
      node234_l = node204_r & ~pixel[241];
      node235_r = node234_l & pixel[528];
      node235_l = node234_l & ~pixel[528];
      node236_r = node235_l & pixel[625];
      node236_l = node235_l & ~pixel[625];
      node237_r = node236_l & pixel[601];
      node237_l = node236_l & ~pixel[601];
      node238 = node237_l;
      node239 = node237_r;
      node240_r = node236_r & pixel[233];
      node240_l = node236_r & ~pixel[233];
      node241 = node240_l;
      node242 = node240_r;
      node243 = node235_r;
      node244_r = node234_r & pixel[371];
      node244_l = node234_r & ~pixel[371];
      node245_r = node244_l & pixel[320];
      node245_l = node244_l & ~pixel[320];
      node246_r = node245_l & pixel[289];
      node246_l = node245_l & ~pixel[289];
      node247 = node246_l;
      node248 = node246_r;
      node249_r = node245_r & pixel[211];
      node249_l = node245_r & ~pixel[211];
      node250 = node249_l;
      node251 = node249_r;
      node252_r = node244_r & pixel[547];
      node252_l = node244_r & ~pixel[547];
      node253_r = node252_l & pixel[262];
      node253_l = node252_l & ~pixel[262];
      node254 = node253_l;
      node255 = node253_r;
      node256_r = node252_r & pixel[267];
      node256_l = node252_r & ~pixel[267];
      node257 = node256_l;
      node258 = node256_r;
      node259_r = node203_r & pixel[344];
      node259_l = node203_r & ~pixel[344];
      node260_r = node259_l & pixel[594];
      node260_l = node259_l & ~pixel[594];
      node261_r = node260_l & pixel[546];
      node261_l = node260_l & ~pixel[546];
      node262_r = node261_l & pixel[398];
      node262_l = node261_l & ~pixel[398];
      node263_r = node262_l & pixel[376];
      node263_l = node262_l & ~pixel[376];
      node264 = node263_l;
      node265 = node263_r;
      node266_r = node262_r & pixel[152];
      node266_l = node262_r & ~pixel[152];
      node267 = node266_l;
      node268 = node266_r;
      node269_r = node261_r & pixel[151];
      node269_l = node261_r & ~pixel[151];
      node270_r = node269_l & pixel[439];
      node270_l = node269_l & ~pixel[439];
      node271 = node270_l;
      node272 = node270_r;
      node273 = node269_r;
      node274_r = node260_r & pixel[493];
      node274_l = node260_r & ~pixel[493];
      node275_r = node274_l & pixel[377];
      node275_l = node274_l & ~pixel[377];
      node276_r = node275_l & pixel[181];
      node276_l = node275_l & ~pixel[181];
      node277 = node276_l;
      node278 = node276_r;
      node279 = node275_r;
      node280_r = node274_r & pixel[377];
      node280_l = node274_r & ~pixel[377];
      node281 = node280_l;
      node282_r = node280_r & pixel[320];
      node282_l = node280_r & ~pixel[320];
      node283 = node282_l;
      node284 = node282_r;
      node285_r = node259_r & pixel[237];
      node285_l = node259_r & ~pixel[237];
      node286_r = node285_l & pixel[411];
      node286_l = node285_l & ~pixel[411];
      node287_r = node286_l & pixel[414];
      node287_l = node286_l & ~pixel[414];
      node288_r = node287_l & pixel[214];
      node288_l = node287_l & ~pixel[214];
      node289 = node288_l;
      node290 = node288_r;
      node291_r = node287_r & pixel[292];
      node291_l = node287_r & ~pixel[292];
      node292 = node291_l;
      node293 = node291_r;
      node294_r = node286_r & pixel[427];
      node294_l = node286_r & ~pixel[427];
      node295_r = node294_l & pixel[576];
      node295_l = node294_l & ~pixel[576];
      node296 = node295_l;
      node297 = node295_r;
      node298_r = node294_r & pixel[360];
      node298_l = node294_r & ~pixel[360];
      node299 = node298_l;
      node300 = node298_r;
      node301_r = node285_r & pixel[215];
      node301_l = node285_r & ~pixel[215];
      node302_r = node301_l & pixel[185];
      node302_l = node301_l & ~pixel[185];
      node303_r = node302_l & pixel[571];
      node303_l = node302_l & ~pixel[571];
      node304 = node303_l;
      node305 = node303_r;
      node306 = node302_r;
      node307_r = node301_r & pixel[240];
      node307_l = node301_r & ~pixel[240];
      node308_r = node307_l & pixel[157];
      node308_l = node307_l & ~pixel[157];
      node309 = node308_l;
      node310 = node308_r;
      node311_r = node307_r & pixel[414];
      node311_l = node307_r & ~pixel[414];
      node312 = node311_l;
      node313 = node311_r;
      node314_r = node202_r & pixel[216];
      node314_l = node202_r & ~pixel[216];
      node315_r = node314_l & pixel[485];
      node315_l = node314_l & ~pixel[485];
      node316_r = node315_l & pixel[275];
      node316_l = node315_l & ~pixel[275];
      node317_r = node316_l & pixel[486];
      node317_l = node316_l & ~pixel[486];
      node318_r = node317_l & pixel[213];
      node318_l = node317_l & ~pixel[213];
      node319_r = node318_l & pixel[179];
      node319_l = node318_l & ~pixel[179];
      node320 = node319_l;
      node321 = node319_r;
      node322_r = node318_r & pixel[348];
      node322_l = node318_r & ~pixel[348];
      node323 = node322_l;
      node324 = node322_r;
      node325_r = node317_r & pixel[243];
      node325_l = node317_r & ~pixel[243];
      node326_r = node325_l & pixel[689];
      node326_l = node325_l & ~pixel[689];
      node327 = node326_l;
      node328 = node326_r;
      node329_r = node325_r & pixel[273];
      node329_l = node325_r & ~pixel[273];
      node330 = node329_l;
      node331 = node329_r;
      node332 = node316_r;
      node333_r = node315_r & pixel[601];
      node333_l = node315_r & ~pixel[601];
      node334_r = node333_l & pixel[376];
      node334_l = node333_l & ~pixel[376];
      node335_r = node334_l & pixel[570];
      node335_l = node334_l & ~pixel[570];
      node336_r = node335_l & pixel[100];
      node336_l = node335_l & ~pixel[100];
      node337 = node336_l;
      node338 = node336_r;
      node339_r = node335_r & pixel[287];
      node339_l = node335_r & ~pixel[287];
      node340 = node339_l;
      node341 = node339_r;
      node342_r = node334_r & pixel[238];
      node342_l = node334_r & ~pixel[238];
      node343 = node342_l;
      node344_r = node342_r & pixel[324];
      node344_l = node342_r & ~pixel[324];
      node345 = node344_l;
      node346 = node344_r;
      node347_r = node333_r & pixel[247];
      node347_l = node333_r & ~pixel[247];
      node348_r = node347_l & pixel[353];
      node348_l = node347_l & ~pixel[353];
      node349_r = node348_l & pixel[164];
      node349_l = node348_l & ~pixel[164];
      node350 = node349_l;
      node351 = node349_r;
      node352_r = node348_r & pixel[234];
      node352_l = node348_r & ~pixel[234];
      node353 = node352_l;
      node354 = node352_r;
      node355_r = node347_r & pixel[397];
      node355_l = node347_r & ~pixel[397];
      node356 = node355_l;
      node357_r = node355_r & pixel[543];
      node357_l = node355_r & ~pixel[543];
      node358 = node357_l;
      node359 = node357_r;
      node360_r = node314_r & pixel[411];
      node360_l = node314_r & ~pixel[411];
      node361_r = node360_l & pixel[517];
      node361_l = node360_l & ~pixel[517];
      node362_r = node361_l & pixel[331];
      node362_l = node361_l & ~pixel[331];
      node363_r = node362_l & pixel[149];
      node363_l = node362_l & ~pixel[149];
      node364_r = node363_l & pixel[127];
      node364_l = node363_l & ~pixel[127];
      node365 = node364_l;
      node366 = node364_r;
      node367_r = node363_r & pixel[400];
      node367_l = node363_r & ~pixel[400];
      node368 = node367_l;
      node369 = node367_r;
      node370_r = node362_r & pixel[385];
      node370_l = node362_r & ~pixel[385];
      node371_r = node370_l & pixel[297];
      node371_l = node370_l & ~pixel[297];
      node372 = node371_l;
      node373 = node371_r;
      node374 = node370_r;
      node375_r = node361_r & pixel[218];
      node375_l = node361_r & ~pixel[218];
      node376_r = node375_l & pixel[212];
      node376_l = node375_l & ~pixel[212];
      node377_r = node376_l & pixel[538];
      node377_l = node376_l & ~pixel[538];
      node378 = node377_l;
      node379 = node377_r;
      node380_r = node376_r & pixel[571];
      node380_l = node376_r & ~pixel[571];
      node381 = node380_l;
      node382 = node380_r;
      node383_r = node375_r & pixel[265];
      node383_l = node375_r & ~pixel[265];
      node384_r = node383_l & pixel[108];
      node384_l = node383_l & ~pixel[108];
      node385 = node384_l;
      node386 = node384_r;
      node387_r = node383_r & pixel[293];
      node387_l = node383_r & ~pixel[293];
      node388 = node387_l;
      node389 = node387_r;
      node390_r = node360_r & pixel[386];
      node390_l = node360_r & ~pixel[386];
      node391_r = node390_l & pixel[657];
      node391_l = node390_l & ~pixel[657];
      node392_r = node391_l & pixel[597];
      node392_l = node391_l & ~pixel[597];
      node393_r = node392_l & pixel[295];
      node393_l = node392_l & ~pixel[295];
      node394 = node393_l;
      node395 = node393_r;
      node396_r = node392_r & pixel[513];
      node396_l = node392_r & ~pixel[513];
      node397 = node396_l;
      node398 = node396_r;
      node399_r = node391_r & pixel[260];
      node399_l = node391_r & ~pixel[260];
      node400_r = node399_l & pixel[238];
      node400_l = node399_l & ~pixel[238];
      node401 = node400_l;
      node402 = node400_r;
      node403 = node399_r;
      node404_r = node390_r & pixel[452];
      node404_l = node390_r & ~pixel[452];
      node405_r = node404_l & pixel[212];
      node405_l = node404_l & ~pixel[212];
      node406 = node405_l;
      node407_r = node405_r & pixel[543];
      node407_l = node405_r & ~pixel[543];
      node408 = node407_l;
      node409 = node407_r;
      node410_r = node404_r & pixel[580];
      node410_l = node404_r & ~pixel[580];
      node411 = node410_l;
      node412 = node410_r;
      node413_r = node1_r & pixel[606];
      node413_l = node1_r & ~pixel[606];
      node414_r = node413_l & pixel[467];
      node414_l = node413_l & ~pixel[467];
      node415_r = node414_l & pixel[318];
      node415_l = node414_l & ~pixel[318];
      node416_r = node415_l & pixel[548];
      node416_l = node415_l & ~pixel[548];
      node417_r = node416_l & pixel[375];
      node417_l = node416_l & ~pixel[375];
      node418_r = node417_l & pixel[714];
      node418_l = node417_l & ~pixel[714];
      node419_r = node418_l & pixel[246];
      node419_l = node418_l & ~pixel[246];
      node420_r = node419_l & pixel[150];
      node420_l = node419_l & ~pixel[150];
      node421 = node420_l;
      node422 = node420_r;
      node423_r = node419_r & pixel[296];
      node423_l = node419_r & ~pixel[296];
      node424 = node423_l;
      node425 = node423_r;
      node426_r = node418_r & pixel[601];
      node426_l = node418_r & ~pixel[601];
      node427_r = node426_l & pixel[377];
      node427_l = node426_l & ~pixel[377];
      node428 = node427_l;
      node429 = node427_r;
      node430_r = node426_r & pixel[352];
      node430_l = node426_r & ~pixel[352];
      node431 = node430_l;
      node432 = node430_r;
      node433_r = node417_r & pixel[183];
      node433_l = node417_r & ~pixel[183];
      node434_r = node433_l & pixel[214];
      node434_l = node433_l & ~pixel[214];
      node435_r = node434_l & pixel[236];
      node435_l = node434_l & ~pixel[236];
      node436 = node435_l;
      node437 = node435_r;
      node438_r = node434_r & pixel[438];
      node438_l = node434_r & ~pixel[438];
      node439 = node438_l;
      node440 = node438_r;
      node441_r = node433_r & pixel[343];
      node441_l = node433_r & ~pixel[343];
      node442_r = node441_l & pixel[516];
      node442_l = node441_l & ~pixel[516];
      node443 = node442_l;
      node444 = node442_r;
      node445_r = node441_r & pixel[517];
      node445_l = node441_r & ~pixel[517];
      node446 = node445_l;
      node447 = node445_r;
      node448_r = node416_r & pixel[521];
      node448_l = node416_r & ~pixel[521];
      node449_r = node448_l & pixel[297];
      node449_l = node448_l & ~pixel[297];
      node450_r = node449_l & pixel[569];
      node450_l = node449_l & ~pixel[569];
      node451_r = node450_l & pixel[659];
      node451_l = node450_l & ~pixel[659];
      node452 = node451_l;
      node453 = node451_r;
      node454_r = node450_r & pixel[461];
      node454_l = node450_r & ~pixel[461];
      node455 = node454_l;
      node456 = node454_r;
      node457_r = node449_r & pixel[271];
      node457_l = node449_r & ~pixel[271];
      node458_r = node457_l & pixel[261];
      node458_l = node457_l & ~pixel[261];
      node459 = node458_l;
      node460 = node458_r;
      node461_r = node457_r & pixel[155];
      node461_l = node457_r & ~pixel[155];
      node462 = node461_l;
      node463 = node461_r;
      node464_r = node448_r & pixel[516];
      node464_l = node448_r & ~pixel[516];
      node465_r = node464_l & pixel[179];
      node465_l = node464_l & ~pixel[179];
      node466_r = node465_l & pixel[626];
      node466_l = node465_l & ~pixel[626];
      node467 = node466_l;
      node468 = node466_r;
      node469_r = node465_r & pixel[293];
      node469_l = node465_r & ~pixel[293];
      node470 = node469_l;
      node471 = node469_r;
      node472_r = node464_r & pixel[524];
      node472_l = node464_r & ~pixel[524];
      node473_r = node472_l & pixel[487];
      node473_l = node472_l & ~pixel[487];
      node474 = node473_l;
      node475 = node473_r;
      node476_r = node472_r & pixel[315];
      node476_l = node472_r & ~pixel[315];
      node477 = node476_l;
      node478 = node476_r;
      node479_r = node415_r & pixel[156];
      node479_l = node415_r & ~pixel[156];
      node480_r = node479_l & pixel[596];
      node480_l = node479_l & ~pixel[596];
      node481_r = node480_l & pixel[577];
      node481_l = node480_l & ~pixel[577];
      node482_r = node481_l & pixel[209];
      node482_l = node481_l & ~pixel[209];
      node483_r = node482_l & pixel[711];
      node483_l = node482_l & ~pixel[711];
      node484 = node483_l;
      node485 = node483_r;
      node486_r = node482_r & pixel[515];
      node486_l = node482_r & ~pixel[515];
      node487 = node486_l;
      node488 = node486_r;
      node489_r = node481_r & pixel[441];
      node489_l = node481_r & ~pixel[441];
      node490_r = node489_l & pixel[657];
      node490_l = node489_l & ~pixel[657];
      node491 = node490_l;
      node492 = node490_r;
      node493_r = node489_r & pixel[321];
      node493_l = node489_r & ~pixel[321];
      node494 = node493_l;
      node495 = node493_r;
      node496_r = node480_r & pixel[681];
      node496_l = node480_r & ~pixel[681];
      node497_r = node496_l & pixel[382];
      node497_l = node496_l & ~pixel[382];
      node498_r = node497_l & pixel[369];
      node498_l = node497_l & ~pixel[369];
      node499 = node498_l;
      node500 = node498_r;
      node501_r = node497_r & pixel[332];
      node501_l = node497_r & ~pixel[332];
      node502 = node501_l;
      node503 = node501_r;
      node504_r = node496_r & pixel[568];
      node504_l = node496_r & ~pixel[568];
      node505_r = node504_l & pixel[326];
      node505_l = node504_l & ~pixel[326];
      node506 = node505_l;
      node507 = node505_r;
      node508_r = node504_r & pixel[486];
      node508_l = node504_r & ~pixel[486];
      node509 = node508_l;
      node510 = node508_r;
      node511_r = node479_r & pixel[458];
      node511_l = node479_r & ~pixel[458];
      node512_r = node511_l & pixel[566];
      node512_l = node511_l & ~pixel[566];
      node513_r = node512_l & pixel[651];
      node513_l = node512_l & ~pixel[651];
      node514_r = node513_l & pixel[571];
      node514_l = node513_l & ~pixel[571];
      node515 = node514_l;
      node516 = node514_r;
      node517_r = node513_r & pixel[274];
      node517_l = node513_r & ~pixel[274];
      node518 = node517_l;
      node519 = node517_r;
      node520_r = node512_r & pixel[440];
      node520_l = node512_r & ~pixel[440];
      node521_r = node520_l & pixel[428];
      node521_l = node520_l & ~pixel[428];
      node522 = node521_l;
      node523 = node521_r;
      node524_r = node520_r & pixel[507];
      node524_l = node520_r & ~pixel[507];
      node525 = node524_l;
      node526 = node524_r;
      node527_r = node511_r & pixel[376];
      node527_l = node511_r & ~pixel[376];
      node528_r = node527_l & pixel[73];
      node528_l = node527_l & ~pixel[73];
      node529_r = node528_l & pixel[463];
      node529_l = node528_l & ~pixel[463];
      node530 = node529_l;
      node531 = node529_r;
      node532 = node528_r;
      node533_r = node527_r & pixel[542];
      node533_l = node527_r & ~pixel[542];
      node534_r = node533_l & pixel[352];
      node534_l = node533_l & ~pixel[352];
      node535 = node534_l;
      node536 = node534_r;
      node537_r = node533_r & pixel[511];
      node537_l = node533_r & ~pixel[511];
      node538 = node537_l;
      node539 = node537_r;
      node540_r = node414_r & pixel[303];
      node540_l = node414_r & ~pixel[303];
      node541_r = node540_l & pixel[527];
      node541_l = node540_l & ~pixel[527];
      node542_r = node541_l & pixel[602];
      node542_l = node541_l & ~pixel[602];
      node543_r = node542_l & pixel[492];
      node543_l = node542_l & ~pixel[492];
      node544_r = node543_l & pixel[523];
      node544_l = node543_l & ~pixel[523];
      node545_r = node544_l & pixel[489];
      node545_l = node544_l & ~pixel[489];
      node546 = node545_l;
      node547 = node545_r;
      node548_r = node544_r & pixel[342];
      node548_l = node544_r & ~pixel[342];
      node549 = node548_l;
      node550 = node548_r;
      node551_r = node543_r & pixel[657];
      node551_l = node543_r & ~pixel[657];
      node552_r = node551_l & pixel[496];
      node552_l = node551_l & ~pixel[496];
      node553 = node552_l;
      node554 = node552_r;
      node555_r = node551_r & pixel[552];
      node555_l = node551_r & ~pixel[552];
      node556 = node555_l;
      node557 = node555_r;
      node558_r = node542_r & pixel[535];
      node558_l = node542_r & ~pixel[535];
      node559_r = node558_l & pixel[516];
      node559_l = node558_l & ~pixel[516];
      node560_r = node559_l & pixel[625];
      node560_l = node559_l & ~pixel[625];
      node561 = node560_l;
      node562 = node560_r;
      node563_r = node559_r & pixel[686];
      node563_l = node559_r & ~pixel[686];
      node564 = node563_l;
      node565 = node563_r;
      node566_r = node558_r & pixel[343];
      node566_l = node558_r & ~pixel[343];
      node567_r = node566_l & pixel[482];
      node567_l = node566_l & ~pixel[482];
      node568 = node567_l;
      node569 = node567_r;
      node570_r = node566_r & pixel[265];
      node570_l = node566_r & ~pixel[265];
      node571 = node570_l;
      node572 = node570_r;
      node573_r = node541_r & pixel[710];
      node573_l = node541_r & ~pixel[710];
      node574_r = node573_l & pixel[355];
      node574_l = node573_l & ~pixel[355];
      node575_r = node574_l & pixel[601];
      node575_l = node574_l & ~pixel[601];
      node576_r = node575_l & pixel[121];
      node576_l = node575_l & ~pixel[121];
      node577 = node576_l;
      node578 = node576_r;
      node579_r = node575_r & pixel[630];
      node579_l = node575_r & ~pixel[630];
      node580 = node579_l;
      node581 = node579_r;
      node582_r = node574_r & pixel[152];
      node582_l = node574_r & ~pixel[152];
      node583_r = node582_l & pixel[176];
      node583_l = node582_l & ~pixel[176];
      node584 = node583_l;
      node585 = node583_r;
      node586_r = node582_r & pixel[381];
      node586_l = node582_r & ~pixel[381];
      node587 = node586_l;
      node588 = node586_r;
      node589 = node573_r;
      node590_r = node540_r & pixel[268];
      node590_l = node540_r & ~pixel[268];
      node591_r = node590_l & pixel[322];
      node591_l = node590_l & ~pixel[322];
      node592_r = node591_l & pixel[352];
      node592_l = node591_l & ~pixel[352];
      node593 = node592_l;
      node594_r = node592_r & pixel[403];
      node594_l = node592_r & ~pixel[403];
      node595 = node594_l;
      node596 = node594_r;
      node597_r = node591_r & pixel[356];
      node597_l = node591_r & ~pixel[356];
      node598 = node597_l;
      node599 = node597_r;
      node600_r = node590_r & pixel[293];
      node600_l = node590_r & ~pixel[293];
      node601_r = node600_l & pixel[372];
      node601_l = node600_l & ~pixel[372];
      node602_r = node601_l & pixel[384];
      node602_l = node601_l & ~pixel[384];
      node603 = node602_l;
      node604 = node602_r;
      node605 = node601_r;
      node606_r = node600_r & pixel[658];
      node606_l = node600_r & ~pixel[658];
      node607 = node606_l;
      node608_r = node606_r & pixel[285];
      node608_l = node606_r & ~pixel[285];
      node609 = node608_l;
      node610 = node608_r;
      node611_r = node413_r & pixel[433];
      node611_l = node413_r & ~pixel[433];
      node612_r = node611_l & pixel[151];
      node612_l = node611_l & ~pixel[151];
      node613_r = node612_l & pixel[245];
      node613_l = node612_l & ~pixel[245];
      node614_r = node613_l & pixel[486];
      node614_l = node613_l & ~pixel[486];
      node615_r = node614_l & pixel[158];
      node615_l = node614_l & ~pixel[158];
      node616_r = node615_l & pixel[600];
      node616_l = node615_l & ~pixel[600];
      node617_r = node616_l & pixel[207];
      node617_l = node616_l & ~pixel[207];
      node618 = node617_l;
      node619 = node617_r;
      node620_r = node616_r & pixel[547];
      node620_l = node616_r & ~pixel[547];
      node621 = node620_l;
      node622 = node620_r;
      node623_r = node615_r & pixel[97];
      node623_l = node615_r & ~pixel[97];
      node624_r = node623_l & pixel[152];
      node624_l = node623_l & ~pixel[152];
      node625 = node624_l;
      node626 = node624_r;
      node627_r = node623_r & pixel[215];
      node627_l = node623_r & ~pixel[215];
      node628 = node627_l;
      node629 = node627_r;
      node630_r = node614_r & pixel[685];
      node630_l = node614_r & ~pixel[685];
      node631_r = node630_l & pixel[572];
      node631_l = node630_l & ~pixel[572];
      node632_r = node631_l & pixel[268];
      node632_l = node631_l & ~pixel[268];
      node633 = node632_l;
      node634 = node632_r;
      node635_r = node631_r & pixel[162];
      node635_l = node631_r & ~pixel[162];
      node636 = node635_l;
      node637 = node635_r;
      node638_r = node630_r & pixel[272];
      node638_l = node630_r & ~pixel[272];
      node639_r = node638_l & pixel[627];
      node639_l = node638_l & ~pixel[627];
      node640 = node639_l;
      node641 = node639_r;
      node642 = node638_r;
      node643_r = node613_r & pixel[458];
      node643_l = node613_r & ~pixel[458];
      node644_r = node643_l & pixel[483];
      node644_l = node643_l & ~pixel[483];
      node645_r = node644_l & pixel[715];
      node645_l = node644_l & ~pixel[715];
      node646_r = node645_l & pixel[301];
      node646_l = node645_l & ~pixel[301];
      node647 = node646_l;
      node648 = node646_r;
      node649 = node645_r;
      node650_r = node644_r & pixel[371];
      node650_l = node644_r & ~pixel[371];
      node651 = node650_l;
      node652_r = node650_r & pixel[238];
      node652_l = node650_r & ~pixel[238];
      node653 = node652_l;
      node654 = node652_r;
      node655_r = node643_r & pixel[401];
      node655_l = node643_r & ~pixel[401];
      node656 = node655_l;
      node657 = node655_r;
      node658_r = node612_r & pixel[458];
      node658_l = node612_r & ~pixel[458];
      node659_r = node658_l & pixel[262];
      node659_l = node658_l & ~pixel[262];
      node660_r = node659_l & pixel[240];
      node660_l = node659_l & ~pixel[240];
      node661_r = node660_l & pixel[343];
      node661_l = node660_l & ~pixel[343];
      node662_r = node661_l & pixel[296];
      node662_l = node661_l & ~pixel[296];
      node663 = node662_l;
      node664 = node662_r;
      node665_r = node661_r & pixel[232];
      node665_l = node661_r & ~pixel[232];
      node666 = node665_l;
      node667 = node665_r;
      node668_r = node660_r & pixel[294];
      node668_l = node660_r & ~pixel[294];
      node669_r = node668_l & pixel[259];
      node669_l = node668_l & ~pixel[259];
      node670 = node669_l;
      node671 = node669_r;
      node672_r = node668_r & pixel[689];
      node672_l = node668_r & ~pixel[689];
      node673 = node672_l;
      node674 = node672_r;
      node675_r = node659_r & pixel[373];
      node675_l = node659_r & ~pixel[373];
      node676_r = node675_l & pixel[270];
      node676_l = node675_l & ~pixel[270];
      node677_r = node676_l & pixel[159];
      node677_l = node676_l & ~pixel[159];
      node678 = node677_l;
      node679 = node677_r;
      node680_r = node676_r & pixel[659];
      node680_l = node676_r & ~pixel[659];
      node681 = node680_l;
      node682 = node680_r;
      node683_r = node675_r & pixel[174];
      node683_l = node675_r & ~pixel[174];
      node684_r = node683_l & pixel[331];
      node684_l = node683_l & ~pixel[331];
      node685 = node684_l;
      node686 = node684_r;
      node687_r = node683_r & pixel[688];
      node687_l = node683_r & ~pixel[688];
      node688 = node687_l;
      node689 = node687_r;
      node690_r = node658_r & pixel[659];
      node690_l = node658_r & ~pixel[659];
      node691_r = node690_l & pixel[328];
      node691_l = node690_l & ~pixel[328];
      node692_r = node691_l & pixel[463];
      node692_l = node691_l & ~pixel[463];
      node693_r = node692_l & pixel[320];
      node693_l = node692_l & ~pixel[320];
      node694 = node693_l;
      node695 = node693_r;
      node696_r = node692_r & pixel[296];
      node696_l = node692_r & ~pixel[296];
      node697 = node696_l;
      node698 = node696_r;
      node699_r = node691_r & pixel[402];
      node699_l = node691_r & ~pixel[402];
      node700 = node699_l;
      node701 = node699_r;
      node702_r = node690_r & pixel[582];
      node702_l = node690_r & ~pixel[582];
      node703_r = node702_l & pixel[489];
      node703_l = node702_l & ~pixel[489];
      node704_r = node703_l & pixel[468];
      node704_l = node703_l & ~pixel[468];
      node705 = node704_l;
      node706 = node704_r;
      node707_r = node703_r & pixel[211];
      node707_l = node703_r & ~pixel[211];
      node708 = node707_l;
      node709 = node707_r;
      node710_r = node702_r & pixel[295];
      node710_l = node702_r & ~pixel[295];
      node711_r = node710_l & pixel[682];
      node711_l = node710_l & ~pixel[682];
      node712 = node711_l;
      node713 = node711_r;
      node714 = node710_r;
      node715_r = node611_r & pixel[610];
      node715_l = node611_r & ~pixel[610];
      node716_r = node715_l & pixel[513];
      node716_l = node715_l & ~pixel[513];
      node717_r = node716_l & pixel[213];
      node717_l = node716_l & ~pixel[213];
      node718_r = node717_l & pixel[261];
      node718_l = node717_l & ~pixel[261];
      node719_r = node718_l & pixel[292];
      node719_l = node718_l & ~pixel[292];
      node720_r = node719_l & pixel[517];
      node720_l = node719_l & ~pixel[517];
      node721 = node720_l;
      node722 = node720_r;
      node723_r = node719_r & pixel[518];
      node723_l = node719_r & ~pixel[518];
      node724 = node723_l;
      node725 = node723_r;
      node726_r = node718_r & pixel[468];
      node726_l = node718_r & ~pixel[468];
      node727_r = node726_l & pixel[547];
      node727_l = node726_l & ~pixel[547];
      node728 = node727_l;
      node729 = node727_r;
      node730_r = node726_r & pixel[583];
      node730_l = node726_r & ~pixel[583];
      node731 = node730_l;
      node732 = node730_r;
      node733_r = node717_r & pixel[517];
      node733_l = node717_r & ~pixel[517];
      node734_r = node733_l & pixel[324];
      node734_l = node733_l & ~pixel[324];
      node735_r = node734_l & pixel[351];
      node735_l = node734_l & ~pixel[351];
      node736 = node735_l;
      node737 = node735_r;
      node738_r = node734_r & pixel[523];
      node738_l = node734_r & ~pixel[523];
      node739 = node738_l;
      node740 = node738_r;
      node741_r = node733_r & pixel[290];
      node741_l = node733_r & ~pixel[290];
      node742_r = node741_l & pixel[347];
      node742_l = node741_l & ~pixel[347];
      node743 = node742_l;
      node744 = node742_r;
      node745_r = node741_r & pixel[581];
      node745_l = node741_r & ~pixel[581];
      node746 = node745_l;
      node747 = node745_r;
      node748_r = node716_r & pixel[384];
      node748_l = node716_r & ~pixel[384];
      node749_r = node748_l & pixel[464];
      node749_l = node748_l & ~pixel[464];
      node750_r = node749_l & pixel[155];
      node750_l = node749_l & ~pixel[155];
      node751_r = node750_l & pixel[359];
      node751_l = node750_l & ~pixel[359];
      node752 = node751_l;
      node753 = node751_r;
      node754_r = node750_r & pixel[291];
      node754_l = node750_r & ~pixel[291];
      node755 = node754_l;
      node756 = node754_r;
      node757_r = node749_r & pixel[298];
      node757_l = node749_r & ~pixel[298];
      node758_r = node757_l & pixel[518];
      node758_l = node757_l & ~pixel[518];
      node759 = node758_l;
      node760 = node758_r;
      node761_r = node757_r & pixel[481];
      node761_l = node757_r & ~pixel[481];
      node762 = node761_l;
      node763 = node761_r;
      node764_r = node748_r & pixel[185];
      node764_l = node748_r & ~pixel[185];
      node765_r = node764_l & pixel[545];
      node765_l = node764_l & ~pixel[545];
      node766_r = node765_l & pixel[570];
      node766_l = node765_l & ~pixel[570];
      node767 = node766_l;
      node768 = node766_r;
      node769 = node765_r;
      node770_r = node764_r & pixel[655];
      node770_l = node764_r & ~pixel[655];
      node771_r = node770_l & pixel[269];
      node771_l = node770_l & ~pixel[269];
      node772 = node771_l;
      node773 = node771_r;
      node774_r = node770_r & pixel[455];
      node774_l = node770_r & ~pixel[455];
      node775 = node774_l;
      node776 = node774_r;
      node777_r = node715_r & pixel[414];
      node777_l = node715_r & ~pixel[414];
      node778_r = node777_l & pixel[346];
      node778_l = node777_l & ~pixel[346];
      node779_r = node778_l & pixel[406];
      node779_l = node778_l & ~pixel[406];
      node780_r = node779_l & pixel[230];
      node780_l = node779_l & ~pixel[230];
      node781_r = node780_l & pixel[657];
      node781_l = node780_l & ~pixel[657];
      node782 = node781_l;
      node783 = node781_r;
      node784_r = node780_r & pixel[210];
      node784_l = node780_r & ~pixel[210];
      node785 = node784_l;
      node786 = node784_r;
      node787_r = node779_r & pixel[372];
      node787_l = node779_r & ~pixel[372];
      node788_r = node787_l & pixel[312];
      node788_l = node787_l & ~pixel[312];
      node789 = node788_l;
      node790 = node788_r;
      node791_r = node787_r & pixel[246];
      node791_l = node787_r & ~pixel[246];
      node792 = node791_l;
      node793 = node791_r;
      node794_r = node778_r & pixel[567];
      node794_l = node778_r & ~pixel[567];
      node795_r = node794_l & pixel[260];
      node795_l = node794_l & ~pixel[260];
      node796_r = node795_l & pixel[572];
      node796_l = node795_l & ~pixel[572];
      node797 = node796_l;
      node798 = node796_r;
      node799_r = node795_r & pixel[557];
      node799_l = node795_r & ~pixel[557];
      node800 = node799_l;
      node801 = node799_r;
      node802 = node794_r;
      node803_r = node777_r & pixel[654];
      node803_l = node777_r & ~pixel[654];
      node804_r = node803_l & pixel[568];
      node804_l = node803_l & ~pixel[568];
      node805_r = node804_l & pixel[574];
      node805_l = node804_l & ~pixel[574];
      node806 = node805_l;
      node807 = node805_r;
      node808_r = node804_r & pixel[328];
      node808_l = node804_r & ~pixel[328];
      node809 = node808_l;
      node810 = node808_r;
      node811_r = node803_r & pixel[429];
      node811_l = node803_r & ~pixel[429];
      node812 = node811_l;
      node813_r = node811_r & pixel[458];
      node813_l = node811_r & ~pixel[458];
      node814 = node813_l;
      node815 = node813_r;
      node816_r = node0_r & pixel[514];
      node816_l = node0_r & ~pixel[514];
      node817_r = node816_l & pixel[157];
      node817_l = node816_l & ~pixel[157];
      node818_r = node817_l & pixel[402];
      node818_l = node817_l & ~pixel[402];
      node819_r = node818_l & pixel[456];
      node819_l = node818_l & ~pixel[456];
      node820_r = node819_l & pixel[405];
      node820_l = node819_l & ~pixel[405];
      node821_r = node820_l & pixel[299];
      node821_l = node820_l & ~pixel[299];
      node822_r = node821_l & pixel[325];
      node822_l = node821_l & ~pixel[325];
      node823_r = node822_l & pixel[709];
      node823_l = node822_l & ~pixel[709];
      node824_r = node823_l & pixel[243];
      node824_l = node823_l & ~pixel[243];
      node825 = node824_l;
      node826 = node824_r;
      node827_r = node823_r & pixel[579];
      node827_l = node823_r & ~pixel[579];
      node828 = node827_l;
      node829 = node827_r;
      node830_r = node822_r & pixel[539];
      node830_l = node822_r & ~pixel[539];
      node831_r = node830_l & pixel[598];
      node831_l = node830_l & ~pixel[598];
      node832 = node831_l;
      node833 = node831_r;
      node834_r = node830_r & pixel[123];
      node834_l = node830_r & ~pixel[123];
      node835 = node834_l;
      node836 = node834_r;
      node837_r = node821_r & pixel[553];
      node837_l = node821_r & ~pixel[553];
      node838_r = node837_l & pixel[154];
      node838_l = node837_l & ~pixel[154];
      node839_r = node838_l & pixel[185];
      node839_l = node838_l & ~pixel[185];
      node840 = node839_l;
      node841 = node839_r;
      node842_r = node838_r & pixel[322];
      node842_l = node838_r & ~pixel[322];
      node843 = node842_l;
      node844 = node842_r;
      node845_r = node837_r & pixel[571];
      node845_l = node837_r & ~pixel[571];
      node846_r = node845_l & pixel[598];
      node846_l = node845_l & ~pixel[598];
      node847 = node846_l;
      node848 = node846_r;
      node849_r = node845_r & pixel[321];
      node849_l = node845_r & ~pixel[321];
      node850 = node849_l;
      node851 = node849_r;
      node852_r = node820_r & pixel[517];
      node852_l = node820_r & ~pixel[517];
      node853_r = node852_l & pixel[177];
      node853_l = node852_l & ~pixel[177];
      node854_r = node853_l & pixel[319];
      node854_l = node853_l & ~pixel[319];
      node855_r = node854_l & pixel[182];
      node855_l = node854_l & ~pixel[182];
      node856 = node855_l;
      node857 = node855_r;
      node858_r = node854_r & pixel[491];
      node858_l = node854_r & ~pixel[491];
      node859 = node858_l;
      node860 = node858_r;
      node861_r = node853_r & pixel[265];
      node861_l = node853_r & ~pixel[265];
      node862_r = node861_l & pixel[290];
      node862_l = node861_l & ~pixel[290];
      node863 = node862_l;
      node864 = node862_r;
      node865_r = node861_r & pixel[272];
      node865_l = node861_r & ~pixel[272];
      node866 = node865_l;
      node867 = node865_r;
      node868_r = node852_r & pixel[154];
      node868_l = node852_r & ~pixel[154];
      node869_r = node868_l & pixel[349];
      node869_l = node868_l & ~pixel[349];
      node870_r = node869_l & pixel[375];
      node870_l = node869_l & ~pixel[375];
      node871 = node870_l;
      node872 = node870_r;
      node873_r = node869_r & pixel[433];
      node873_l = node869_r & ~pixel[433];
      node874 = node873_l;
      node875 = node873_r;
      node876_r = node868_r & pixel[178];
      node876_l = node868_r & ~pixel[178];
      node877_r = node876_l & pixel[573];
      node877_l = node876_l & ~pixel[573];
      node878 = node877_l;
      node879 = node877_r;
      node880_r = node876_r & pixel[375];
      node880_l = node876_r & ~pixel[375];
      node881 = node880_l;
      node882 = node880_r;
      node883_r = node819_r & pixel[457];
      node883_l = node819_r & ~pixel[457];
      node884_r = node883_l & pixel[70];
      node884_l = node883_l & ~pixel[70];
      node885_r = node884_l & pixel[597];
      node885_l = node884_l & ~pixel[597];
      node886_r = node885_l & pixel[652];
      node886_l = node885_l & ~pixel[652];
      node887 = node886_l;
      node888 = node886_r;
      node889_r = node885_r & pixel[295];
      node889_l = node885_r & ~pixel[295];
      node890_r = node889_l & pixel[377];
      node890_l = node889_l & ~pixel[377];
      node891 = node890_l;
      node892 = node890_r;
      node893_r = node889_r & pixel[609];
      node893_l = node889_r & ~pixel[609];
      node894 = node893_l;
      node895 = node893_r;
      node896 = node884_r;
      node897_r = node883_r & pixel[264];
      node897_l = node883_r & ~pixel[264];
      node898_r = node897_l & pixel[182];
      node898_l = node897_l & ~pixel[182];
      node899_r = node898_l & pixel[238];
      node899_l = node898_l & ~pixel[238];
      node900_r = node899_l & pixel[123];
      node900_l = node899_l & ~pixel[123];
      node901 = node900_l;
      node902 = node900_r;
      node903_r = node899_r & pixel[484];
      node903_l = node899_r & ~pixel[484];
      node904 = node903_l;
      node905 = node903_r;
      node906_r = node898_r & pixel[371];
      node906_l = node898_r & ~pixel[371];
      node907_r = node906_l & pixel[512];
      node907_l = node906_l & ~pixel[512];
      node908 = node907_l;
      node909 = node907_r;
      node910_r = node906_r & pixel[185];
      node910_l = node906_r & ~pixel[185];
      node911 = node910_l;
      node912 = node910_r;
      node913_r = node897_r & pixel[537];
      node913_l = node897_r & ~pixel[537];
      node914_r = node913_l & pixel[212];
      node914_l = node913_l & ~pixel[212];
      node915_r = node914_l & pixel[217];
      node915_l = node914_l & ~pixel[217];
      node916 = node915_l;
      node917 = node915_r;
      node918_r = node914_r & pixel[299];
      node918_l = node914_r & ~pixel[299];
      node919 = node918_l;
      node920 = node918_r;
      node921_r = node913_r & pixel[238];
      node921_l = node913_r & ~pixel[238];
      node922_r = node921_l & pixel[688];
      node922_l = node921_l & ~pixel[688];
      node923 = node922_l;
      node924 = node922_r;
      node925_r = node921_r & pixel[715];
      node925_l = node921_r & ~pixel[715];
      node926 = node925_l;
      node927 = node925_r;
      node928_r = node818_r & pixel[211];
      node928_l = node818_r & ~pixel[211];
      node929_r = node928_l & pixel[624];
      node929_l = node928_l & ~pixel[624];
      node930_r = node929_l & pixel[433];
      node930_l = node929_l & ~pixel[433];
      node931_r = node930_l & pixel[293];
      node931_l = node930_l & ~pixel[293];
      node932_r = node931_l & pixel[742];
      node932_l = node931_l & ~pixel[742];
      node933_r = node932_l & pixel[127];
      node933_l = node932_l & ~pixel[127];
      node934 = node933_l;
      node935 = node933_r;
      node936_r = node932_r & pixel[351];
      node936_l = node932_r & ~pixel[351];
      node937 = node936_l;
      node938 = node936_r;
      node939_r = node931_r & pixel[317];
      node939_l = node931_r & ~pixel[317];
      node940_r = node939_l & pixel[567];
      node940_l = node939_l & ~pixel[567];
      node941 = node940_l;
      node942 = node940_r;
      node943_r = node939_r & pixel[268];
      node943_l = node939_r & ~pixel[268];
      node944 = node943_l;
      node945 = node943_r;
      node946_r = node930_r & pixel[743];
      node946_l = node930_r & ~pixel[743];
      node947_r = node946_l & pixel[295];
      node947_l = node946_l & ~pixel[295];
      node948_r = node947_l & pixel[491];
      node948_l = node947_l & ~pixel[491];
      node949 = node948_l;
      node950 = node948_r;
      node951_r = node947_r & pixel[523];
      node951_l = node947_r & ~pixel[523];
      node952 = node951_l;
      node953 = node951_r;
      node954_r = node946_r & pixel[521];
      node954_l = node946_r & ~pixel[521];
      node955_r = node954_l & pixel[742];
      node955_l = node954_l & ~pixel[742];
      node956 = node955_l;
      node957 = node955_r;
      node958_r = node954_r & pixel[257];
      node958_l = node954_r & ~pixel[257];
      node959 = node958_l;
      node960 = node958_r;
      node961_r = node929_r & pixel[353];
      node961_l = node929_r & ~pixel[353];
      node962_r = node961_l & pixel[357];
      node962_l = node961_l & ~pixel[357];
      node963_r = node962_l & pixel[180];
      node963_l = node962_l & ~pixel[180];
      node964_r = node963_l & pixel[136];
      node964_l = node963_l & ~pixel[136];
      node965 = node964_l;
      node966 = node964_r;
      node967 = node963_r;
      node968_r = node962_r & pixel[193];
      node968_l = node962_r & ~pixel[193];
      node969_r = node968_l & pixel[360];
      node969_l = node968_l & ~pixel[360];
      node970 = node969_l;
      node971 = node969_r;
      node972 = node968_r;
      node973_r = node961_r & pixel[323];
      node973_l = node961_r & ~pixel[323];
      node974_r = node973_l & pixel[102];
      node974_l = node973_l & ~pixel[102];
      node975_r = node974_l & pixel[553];
      node975_l = node974_l & ~pixel[553];
      node976 = node975_l;
      node977 = node975_r;
      node978 = node974_r;
      node979_r = node973_r & pixel[602];
      node979_l = node973_r & ~pixel[602];
      node980_r = node979_l & pixel[432];
      node980_l = node979_l & ~pixel[432];
      node981 = node980_l;
      node982 = node980_r;
      node983_r = node979_r & pixel[594];
      node983_l = node979_r & ~pixel[594];
      node984 = node983_l;
      node985 = node983_r;
      node986_r = node928_r & pixel[317];
      node986_l = node928_r & ~pixel[317];
      node987_r = node986_l & pixel[349];
      node987_l = node986_l & ~pixel[349];
      node988_r = node987_l & pixel[595];
      node988_l = node987_l & ~pixel[595];
      node989_r = node988_l & pixel[511];
      node989_l = node988_l & ~pixel[511];
      node990_r = node989_l & pixel[208];
      node990_l = node989_l & ~pixel[208];
      node991 = node990_l;
      node992 = node990_r;
      node993_r = node989_r & pixel[377];
      node993_l = node989_r & ~pixel[377];
      node994 = node993_l;
      node995 = node993_r;
      node996_r = node988_r & pixel[555];
      node996_l = node988_r & ~pixel[555];
      node997_r = node996_l & pixel[297];
      node997_l = node996_l & ~pixel[297];
      node998 = node997_l;
      node999 = node997_r;
      node1000_r = node996_r & pixel[343];
      node1000_l = node996_r & ~pixel[343];
      node1001 = node1000_l;
      node1002 = node1000_r;
      node1003_r = node987_r & pixel[190];
      node1003_l = node987_r & ~pixel[190];
      node1004_r = node1003_l & pixel[177];
      node1004_l = node1003_l & ~pixel[177];
      node1005_r = node1004_l & pixel[464];
      node1005_l = node1004_l & ~pixel[464];
      node1006 = node1005_l;
      node1007 = node1005_r;
      node1008_r = node1004_r & pixel[693];
      node1008_l = node1004_r & ~pixel[693];
      node1009 = node1008_l;
      node1010 = node1008_r;
      node1011_r = node1003_r & pixel[484];
      node1011_l = node1003_r & ~pixel[484];
      node1012_r = node1011_l & pixel[324];
      node1012_l = node1011_l & ~pixel[324];
      node1013 = node1012_l;
      node1014 = node1012_r;
      node1015_r = node1011_r & pixel[215];
      node1015_l = node1011_r & ~pixel[215];
      node1016 = node1015_l;
      node1017 = node1015_r;
      node1018_r = node986_r & pixel[191];
      node1018_l = node986_r & ~pixel[191];
      node1019_r = node1018_l & pixel[470];
      node1019_l = node1018_l & ~pixel[470];
      node1020_r = node1019_l & pixel[153];
      node1020_l = node1019_l & ~pixel[153];
      node1021_r = node1020_l & pixel[325];
      node1021_l = node1020_l & ~pixel[325];
      node1022 = node1021_l;
      node1023 = node1021_r;
      node1024_r = node1020_r & pixel[630];
      node1024_l = node1020_r & ~pixel[630];
      node1025 = node1024_l;
      node1026 = node1024_r;
      node1027_r = node1019_r & pixel[206];
      node1027_l = node1019_r & ~pixel[206];
      node1028_r = node1027_l & pixel[119];
      node1028_l = node1027_l & ~pixel[119];
      node1029 = node1028_l;
      node1030 = node1028_r;
      node1031_r = node1027_r & pixel[293];
      node1031_l = node1027_r & ~pixel[293];
      node1032 = node1031_l;
      node1033 = node1031_r;
      node1034_r = node1018_r & pixel[385];
      node1034_l = node1018_r & ~pixel[385];
      node1035_r = node1034_l & pixel[603];
      node1035_l = node1034_l & ~pixel[603];
      node1036_r = node1035_l & pixel[299];
      node1036_l = node1035_l & ~pixel[299];
      node1037 = node1036_l;
      node1038 = node1036_r;
      node1039_r = node1035_r & pixel[188];
      node1039_l = node1035_r & ~pixel[188];
      node1040 = node1039_l;
      node1041 = node1039_r;
      node1042_r = node1034_r & pixel[551];
      node1042_l = node1034_r & ~pixel[551];
      node1043_r = node1042_l & pixel[537];
      node1043_l = node1042_l & ~pixel[537];
      node1044 = node1043_l;
      node1045 = node1043_r;
      node1046_r = node1042_r & pixel[299];
      node1046_l = node1042_r & ~pixel[299];
      node1047 = node1046_l;
      node1048 = node1046_r;
      node1049_r = node817_r & pixel[324];
      node1049_l = node817_r & ~pixel[324];
      node1050_r = node1049_l & pixel[518];
      node1050_l = node1049_l & ~pixel[518];
      node1051_r = node1050_l & pixel[290];
      node1051_l = node1050_l & ~pixel[290];
      node1052_r = node1051_l & pixel[241];
      node1052_l = node1051_l & ~pixel[241];
      node1053_r = node1052_l & pixel[329];
      node1053_l = node1052_l & ~pixel[329];
      node1054_r = node1053_l & pixel[272];
      node1054_l = node1053_l & ~pixel[272];
      node1055_r = node1054_l & pixel[515];
      node1055_l = node1054_l & ~pixel[515];
      node1056 = node1055_l;
      node1057 = node1055_r;
      node1058_r = node1054_r & pixel[380];
      node1058_l = node1054_r & ~pixel[380];
      node1059 = node1058_l;
      node1060 = node1058_r;
      node1061_r = node1053_r & pixel[516];
      node1061_l = node1053_r & ~pixel[516];
      node1062_r = node1061_l & pixel[483];
      node1062_l = node1061_l & ~pixel[483];
      node1063 = node1062_l;
      node1064 = node1062_r;
      node1065 = node1061_r;
      node1066_r = node1052_r & pixel[380];
      node1066_l = node1052_r & ~pixel[380];
      node1067_r = node1066_l & pixel[343];
      node1067_l = node1066_l & ~pixel[343];
      node1068_r = node1067_l & pixel[599];
      node1068_l = node1067_l & ~pixel[599];
      node1069 = node1068_l;
      node1070 = node1068_r;
      node1071 = node1067_r;
      node1072_r = node1066_r & pixel[314];
      node1072_l = node1066_r & ~pixel[314];
      node1073_r = node1072_l & pixel[484];
      node1073_l = node1072_l & ~pixel[484];
      node1074 = node1073_l;
      node1075 = node1073_r;
      node1076_r = node1072_r & pixel[624];
      node1076_l = node1072_r & ~pixel[624];
      node1077 = node1076_l;
      node1078 = node1076_r;
      node1079_r = node1051_r & pixel[457];
      node1079_l = node1051_r & ~pixel[457];
      node1080_r = node1079_l & pixel[301];
      node1080_l = node1079_l & ~pixel[301];
      node1081_r = node1080_l & pixel[211];
      node1081_l = node1080_l & ~pixel[211];
      node1082_r = node1081_l & pixel[267];
      node1082_l = node1081_l & ~pixel[267];
      node1083 = node1082_l;
      node1084 = node1082_r;
      node1085_r = node1081_r & pixel[499];
      node1085_l = node1081_r & ~pixel[499];
      node1086 = node1085_l;
      node1087 = node1085_r;
      node1088_r = node1080_r & pixel[380];
      node1088_l = node1080_r & ~pixel[380];
      node1089 = node1088_l;
      node1090_r = node1088_r & pixel[372];
      node1090_l = node1088_r & ~pixel[372];
      node1091 = node1090_l;
      node1092 = node1090_r;
      node1093_r = node1079_r & pixel[540];
      node1093_l = node1079_r & ~pixel[540];
      node1094_r = node1093_l & pixel[481];
      node1094_l = node1093_l & ~pixel[481];
      node1095_r = node1094_l & pixel[328];
      node1095_l = node1094_l & ~pixel[328];
      node1096 = node1095_l;
      node1097 = node1095_r;
      node1098_r = node1094_r & pixel[302];
      node1098_l = node1094_r & ~pixel[302];
      node1099 = node1098_l;
      node1100 = node1098_r;
      node1101_r = node1093_r & pixel[469];
      node1101_l = node1093_r & ~pixel[469];
      node1102_r = node1101_l & pixel[269];
      node1102_l = node1101_l & ~pixel[269];
      node1103 = node1102_l;
      node1104 = node1102_r;
      node1105_r = node1101_r & pixel[655];
      node1105_l = node1101_r & ~pixel[655];
      node1106 = node1105_l;
      node1107 = node1105_r;
      node1108_r = node1050_r & pixel[349];
      node1108_l = node1050_r & ~pixel[349];
      node1109_r = node1108_l & pixel[566];
      node1109_l = node1108_l & ~pixel[566];
      node1110_r = node1109_l & pixel[345];
      node1110_l = node1109_l & ~pixel[345];
      node1111_r = node1110_l & pixel[264];
      node1111_l = node1110_l & ~pixel[264];
      node1112_r = node1111_l & pixel[689];
      node1112_l = node1111_l & ~pixel[689];
      node1113 = node1112_l;
      node1114 = node1112_r;
      node1115_r = node1111_r & pixel[468];
      node1115_l = node1111_r & ~pixel[468];
      node1116 = node1115_l;
      node1117 = node1115_r;
      node1118_r = node1110_r & pixel[686];
      node1118_l = node1110_r & ~pixel[686];
      node1119_r = node1118_l & pixel[540];
      node1119_l = node1118_l & ~pixel[540];
      node1120 = node1119_l;
      node1121 = node1119_r;
      node1122_r = node1118_r & pixel[485];
      node1122_l = node1118_r & ~pixel[485];
      node1123 = node1122_l;
      node1124 = node1122_r;
      node1125_r = node1109_r & pixel[348];
      node1125_l = node1109_r & ~pixel[348];
      node1126_r = node1125_l & pixel[432];
      node1126_l = node1125_l & ~pixel[432];
      node1127_r = node1126_l & pixel[292];
      node1127_l = node1126_l & ~pixel[292];
      node1128 = node1127_l;
      node1129 = node1127_r;
      node1130_r = node1126_r & pixel[602];
      node1130_l = node1126_r & ~pixel[602];
      node1131 = node1130_l;
      node1132 = node1130_r;
      node1133_r = node1125_r & pixel[433];
      node1133_l = node1125_r & ~pixel[433];
      node1134_r = node1133_l & pixel[627];
      node1134_l = node1133_l & ~pixel[627];
      node1135 = node1134_l;
      node1136 = node1134_r;
      node1137_r = node1133_r & pixel[488];
      node1137_l = node1133_r & ~pixel[488];
      node1138 = node1137_l;
      node1139 = node1137_r;
      node1140_r = node1108_r & pixel[405];
      node1140_l = node1108_r & ~pixel[405];
      node1141_r = node1140_l & pixel[243];
      node1141_l = node1140_l & ~pixel[243];
      node1142_r = node1141_l & pixel[218];
      node1142_l = node1141_l & ~pixel[218];
      node1143_r = node1142_l & pixel[478];
      node1143_l = node1142_l & ~pixel[478];
      node1144 = node1143_l;
      node1145 = node1143_r;
      node1146_r = node1142_r & pixel[461];
      node1146_l = node1142_r & ~pixel[461];
      node1147 = node1146_l;
      node1148 = node1146_r;
      node1149_r = node1141_r & pixel[403];
      node1149_l = node1141_r & ~pixel[403];
      node1150_r = node1149_l & pixel[520];
      node1150_l = node1149_l & ~pixel[520];
      node1151 = node1150_l;
      node1152 = node1150_r;
      node1153_r = node1149_r & pixel[455];
      node1153_l = node1149_r & ~pixel[455];
      node1154 = node1153_l;
      node1155 = node1153_r;
      node1156_r = node1140_r & pixel[355];
      node1156_l = node1140_r & ~pixel[355];
      node1157_r = node1156_l & pixel[263];
      node1157_l = node1156_l & ~pixel[263];
      node1158_r = node1157_l & pixel[235];
      node1158_l = node1157_l & ~pixel[235];
      node1159 = node1158_l;
      node1160 = node1158_r;
      node1161_r = node1157_r & pixel[597];
      node1161_l = node1157_r & ~pixel[597];
      node1162 = node1161_l;
      node1163 = node1161_r;
      node1164_r = node1156_r & pixel[482];
      node1164_l = node1156_r & ~pixel[482];
      node1165_r = node1164_l & pixel[630];
      node1165_l = node1164_l & ~pixel[630];
      node1166 = node1165_l;
      node1167 = node1165_r;
      node1168_r = node1164_r & pixel[320];
      node1168_l = node1164_r & ~pixel[320];
      node1169 = node1168_l;
      node1170 = node1168_r;
      node1171_r = node1049_r & pixel[626];
      node1171_l = node1049_r & ~pixel[626];
      node1172_r = node1171_l & pixel[650];
      node1172_l = node1171_l & ~pixel[650];
      node1173_r = node1172_l & pixel[682];
      node1173_l = node1172_l & ~pixel[682];
      node1174_r = node1173_l & pixel[627];
      node1174_l = node1173_l & ~pixel[627];
      node1175_r = node1174_l & pixel[268];
      node1175_l = node1174_l & ~pixel[268];
      node1176_r = node1175_l & pixel[571];
      node1176_l = node1175_l & ~pixel[571];
      node1177 = node1176_l;
      node1178 = node1176_r;
      node1179_r = node1175_r & pixel[600];
      node1179_l = node1175_r & ~pixel[600];
      node1180 = node1179_l;
      node1181 = node1179_r;
      node1182_r = node1174_r & pixel[634];
      node1182_l = node1174_r & ~pixel[634];
      node1183_r = node1182_l & pixel[346];
      node1183_l = node1182_l & ~pixel[346];
      node1184 = node1183_l;
      node1185 = node1183_r;
      node1186_r = node1182_r & pixel[293];
      node1186_l = node1182_r & ~pixel[293];
      node1187 = node1186_l;
      node1188 = node1186_r;
      node1189_r = node1173_r & pixel[238];
      node1189_l = node1173_r & ~pixel[238];
      node1190_r = node1189_l & pixel[629];
      node1190_l = node1189_l & ~pixel[629];
      node1191_r = node1190_l & pixel[583];
      node1191_l = node1190_l & ~pixel[583];
      node1192 = node1191_l;
      node1193 = node1191_r;
      node1194_r = node1190_r & pixel[685];
      node1194_l = node1190_r & ~pixel[685];
      node1195 = node1194_l;
      node1196 = node1194_r;
      node1197_r = node1189_r & pixel[353];
      node1197_l = node1189_r & ~pixel[353];
      node1198 = node1197_l;
      node1199 = node1197_r;
      node1200_r = node1172_r & pixel[292];
      node1200_l = node1172_r & ~pixel[292];
      node1201_r = node1200_l & pixel[190];
      node1201_l = node1200_l & ~pixel[190];
      node1202 = node1201_l;
      node1203_r = node1201_r & pixel[317];
      node1203_l = node1201_r & ~pixel[317];
      node1204 = node1203_l;
      node1205 = node1203_r;
      node1206_r = node1200_r & pixel[686];
      node1206_l = node1200_r & ~pixel[686];
      node1207 = node1206_l;
      node1208_r = node1206_r & pixel[151];
      node1208_l = node1206_r & ~pixel[151];
      node1209_r = node1208_l & pixel[351];
      node1209_l = node1208_l & ~pixel[351];
      node1210 = node1209_l;
      node1211 = node1209_r;
      node1212 = node1208_r;
      node1213_r = node1171_r & pixel[516];
      node1213_l = node1171_r & ~pixel[516];
      node1214_r = node1213_l & pixel[263];
      node1214_l = node1213_l & ~pixel[263];
      node1215_r = node1214_l & pixel[259];
      node1215_l = node1214_l & ~pixel[259];
      node1216_r = node1215_l & pixel[406];
      node1216_l = node1215_l & ~pixel[406];
      node1217_r = node1216_l & pixel[154];
      node1217_l = node1216_l & ~pixel[154];
      node1218 = node1217_l;
      node1219 = node1217_r;
      node1220_r = node1216_r & pixel[150];
      node1220_l = node1216_r & ~pixel[150];
      node1221 = node1220_l;
      node1222 = node1220_r;
      node1223_r = node1215_r & pixel[346];
      node1223_l = node1215_r & ~pixel[346];
      node1224_r = node1223_l & pixel[350];
      node1224_l = node1223_l & ~pixel[350];
      node1225 = node1224_l;
      node1226 = node1224_r;
      node1227_r = node1223_r & pixel[242];
      node1227_l = node1223_r & ~pixel[242];
      node1228 = node1227_l;
      node1229 = node1227_r;
      node1230_r = node1214_r & pixel[432];
      node1230_l = node1214_r & ~pixel[432];
      node1231_r = node1230_l & pixel[271];
      node1231_l = node1230_l & ~pixel[271];
      node1232_r = node1231_l & pixel[520];
      node1232_l = node1231_l & ~pixel[520];
      node1233 = node1232_l;
      node1234 = node1232_r;
      node1235_r = node1231_r & pixel[345];
      node1235_l = node1231_r & ~pixel[345];
      node1236 = node1235_l;
      node1237 = node1235_r;
      node1238_r = node1230_r & pixel[319];
      node1238_l = node1230_r & ~pixel[319];
      node1239_r = node1238_l & pixel[683];
      node1239_l = node1238_l & ~pixel[683];
      node1240 = node1239_l;
      node1241 = node1239_r;
      node1242_r = node1238_r & pixel[270];
      node1242_l = node1238_r & ~pixel[270];
      node1243 = node1242_l;
      node1244 = node1242_r;
      node1245_r = node1213_r & pixel[569];
      node1245_l = node1213_r & ~pixel[569];
      node1246_r = node1245_l & pixel[604];
      node1246_l = node1245_l & ~pixel[604];
      node1247_r = node1246_l & pixel[180];
      node1247_l = node1246_l & ~pixel[180];
      node1248_r = node1247_l & pixel[292];
      node1248_l = node1247_l & ~pixel[292];
      node1249 = node1248_l;
      node1250 = node1248_r;
      node1251_r = node1247_r & pixel[406];
      node1251_l = node1247_r & ~pixel[406];
      node1252 = node1251_l;
      node1253 = node1251_r;
      node1254_r = node1246_r & pixel[147];
      node1254_l = node1246_r & ~pixel[147];
      node1255_r = node1254_l & pixel[149];
      node1255_l = node1254_l & ~pixel[149];
      node1256 = node1255_l;
      node1257 = node1255_r;
      node1258 = node1254_r;
      node1259_r = node1245_r & pixel[127];
      node1259_l = node1245_r & ~pixel[127];
      node1260_r = node1259_l & pixel[210];
      node1260_l = node1259_l & ~pixel[210];
      node1261_r = node1260_l & pixel[272];
      node1261_l = node1260_l & ~pixel[272];
      node1262 = node1261_l;
      node1263 = node1261_r;
      node1264_r = node1260_r & pixel[574];
      node1264_l = node1260_r & ~pixel[574];
      node1265 = node1264_l;
      node1266 = node1264_r;
      node1267_r = node1259_r & pixel[376];
      node1267_l = node1259_r & ~pixel[376];
      node1268_r = node1267_l & pixel[297];
      node1268_l = node1267_l & ~pixel[297];
      node1269 = node1268_l;
      node1270 = node1268_r;
      node1271_r = node1267_r & pixel[293];
      node1271_l = node1267_r & ~pixel[293];
      node1272 = node1271_l;
      node1273 = node1271_r;
      node1274_r = node816_r & pixel[101];
      node1274_l = node816_r & ~pixel[101];
      node1275_r = node1274_l & pixel[683];
      node1275_l = node1274_l & ~pixel[683];
      node1276_r = node1275_l & pixel[97];
      node1276_l = node1275_l & ~pixel[97];
      node1277_r = node1276_l & pixel[371];
      node1277_l = node1276_l & ~pixel[371];
      node1278_r = node1277_l & pixel[347];
      node1278_l = node1277_l & ~pixel[347];
      node1279_r = node1278_l & pixel[350];
      node1279_l = node1278_l & ~pixel[350];
      node1280_r = node1279_l & pixel[680];
      node1280_l = node1279_l & ~pixel[680];
      node1281_r = node1280_l & pixel[188];
      node1281_l = node1280_l & ~pixel[188];
      node1282 = node1281_l;
      node1283 = node1281_r;
      node1284_r = node1280_r & pixel[155];
      node1284_l = node1280_r & ~pixel[155];
      node1285 = node1284_l;
      node1286 = node1284_r;
      node1287_r = node1279_r & pixel[154];
      node1287_l = node1279_r & ~pixel[154];
      node1288_r = node1287_l & pixel[465];
      node1288_l = node1287_l & ~pixel[465];
      node1289 = node1288_l;
      node1290 = node1288_r;
      node1291_r = node1287_r & pixel[205];
      node1291_l = node1287_r & ~pixel[205];
      node1292 = node1291_l;
      node1293 = node1291_r;
      node1294_r = node1278_r & pixel[405];
      node1294_l = node1278_r & ~pixel[405];
      node1295_r = node1294_l & pixel[655];
      node1295_l = node1294_l & ~pixel[655];
      node1296_r = node1295_l & pixel[600];
      node1296_l = node1295_l & ~pixel[600];
      node1297 = node1296_l;
      node1298 = node1296_r;
      node1299_r = node1295_r & pixel[490];
      node1299_l = node1295_r & ~pixel[490];
      node1300 = node1299_l;
      node1301 = node1299_r;
      node1302_r = node1294_r & pixel[374];
      node1302_l = node1294_r & ~pixel[374];
      node1303_r = node1302_l & pixel[627];
      node1303_l = node1302_l & ~pixel[627];
      node1304 = node1303_l;
      node1305 = node1303_r;
      node1306_r = node1302_r & pixel[271];
      node1306_l = node1302_r & ~pixel[271];
      node1307 = node1306_l;
      node1308 = node1306_r;
      node1309_r = node1277_r & pixel[242];
      node1309_l = node1277_r & ~pixel[242];
      node1310_r = node1309_l & pixel[246];
      node1310_l = node1309_l & ~pixel[246];
      node1311_r = node1310_l & pixel[414];
      node1311_l = node1310_l & ~pixel[414];
      node1312_r = node1311_l & pixel[601];
      node1312_l = node1311_l & ~pixel[601];
      node1313 = node1312_l;
      node1314 = node1312_r;
      node1315_r = node1311_r & pixel[549];
      node1315_l = node1311_r & ~pixel[549];
      node1316 = node1315_l;
      node1317 = node1315_r;
      node1318_r = node1310_r & pixel[183];
      node1318_l = node1310_r & ~pixel[183];
      node1319_r = node1318_l & pixel[217];
      node1319_l = node1318_l & ~pixel[217];
      node1320 = node1319_l;
      node1321 = node1319_r;
      node1322_r = node1318_r & pixel[425];
      node1322_l = node1318_r & ~pixel[425];
      node1323 = node1322_l;
      node1324 = node1322_r;
      node1325_r = node1309_r & pixel[718];
      node1325_l = node1309_r & ~pixel[718];
      node1326_r = node1325_l & pixel[599];
      node1326_l = node1325_l & ~pixel[599];
      node1327_r = node1326_l & pixel[686];
      node1327_l = node1326_l & ~pixel[686];
      node1328 = node1327_l;
      node1329 = node1327_r;
      node1330_r = node1326_r & pixel[405];
      node1330_l = node1326_r & ~pixel[405];
      node1331 = node1330_l;
      node1332 = node1330_r;
      node1333_r = node1325_r & pixel[183];
      node1333_l = node1325_r & ~pixel[183];
      node1334_r = node1333_l & pixel[239];
      node1334_l = node1333_l & ~pixel[239];
      node1335 = node1334_l;
      node1336 = node1334_r;
      node1337_r = node1333_r & pixel[526];
      node1337_l = node1333_r & ~pixel[526];
      node1338 = node1337_l;
      node1339 = node1337_r;
      node1340_r = node1276_r & pixel[440];
      node1340_l = node1276_r & ~pixel[440];
      node1341_r = node1340_l & pixel[415];
      node1341_l = node1340_l & ~pixel[415];
      node1342_r = node1341_l & pixel[291];
      node1342_l = node1341_l & ~pixel[291];
      node1343_r = node1342_l & pixel[386];
      node1343_l = node1342_l & ~pixel[386];
      node1344_r = node1343_l & pixel[517];
      node1344_l = node1343_l & ~pixel[517];
      node1345 = node1344_l;
      node1346 = node1344_r;
      node1347 = node1343_r;
      node1348_r = node1342_r & pixel[297];
      node1348_l = node1342_r & ~pixel[297];
      node1349_r = node1348_l & pixel[607];
      node1349_l = node1348_l & ~pixel[607];
      node1350 = node1349_l;
      node1351 = node1349_r;
      node1352_r = node1348_r & pixel[156];
      node1352_l = node1348_r & ~pixel[156];
      node1353 = node1352_l;
      node1354 = node1352_r;
      node1355_r = node1341_r & pixel[357];
      node1355_l = node1341_r & ~pixel[357];
      node1356_r = node1355_l & pixel[517];
      node1356_l = node1355_l & ~pixel[517];
      node1357 = node1356_l;
      node1358 = node1356_r;
      node1359 = node1355_r;
      node1360_r = node1340_r & pixel[510];
      node1360_l = node1340_r & ~pixel[510];
      node1361_r = node1360_l & pixel[595];
      node1361_l = node1360_l & ~pixel[595];
      node1362_r = node1361_l & pixel[157];
      node1362_l = node1361_l & ~pixel[157];
      node1363_r = node1362_l & pixel[270];
      node1363_l = node1362_l & ~pixel[270];
      node1364 = node1363_l;
      node1365 = node1363_r;
      node1366_r = node1362_r & pixel[317];
      node1366_l = node1362_r & ~pixel[317];
      node1367 = node1366_l;
      node1368 = node1366_r;
      node1369_r = node1361_r & pixel[605];
      node1369_l = node1361_r & ~pixel[605];
      node1370_r = node1369_l & pixel[631];
      node1370_l = node1369_l & ~pixel[631];
      node1371 = node1370_l;
      node1372 = node1370_r;
      node1373 = node1369_r;
      node1374_r = node1360_r & pixel[413];
      node1374_l = node1360_r & ~pixel[413];
      node1375_r = node1374_l & pixel[320];
      node1375_l = node1374_l & ~pixel[320];
      node1376 = node1375_l;
      node1377_r = node1375_r & pixel[343];
      node1377_l = node1375_r & ~pixel[343];
      node1378 = node1377_l;
      node1379 = node1377_r;
      node1380_r = node1374_r & pixel[213];
      node1380_l = node1374_r & ~pixel[213];
      node1381_r = node1380_l & pixel[207];
      node1381_l = node1380_l & ~pixel[207];
      node1382 = node1381_l;
      node1383 = node1381_r;
      node1384_r = node1380_r & pixel[352];
      node1384_l = node1380_r & ~pixel[352];
      node1385 = node1384_l;
      node1386 = node1384_r;
      node1387_r = node1275_r & pixel[541];
      node1387_l = node1275_r & ~pixel[541];
      node1388_r = node1387_l & pixel[212];
      node1388_l = node1387_l & ~pixel[212];
      node1389_r = node1388_l & pixel[600];
      node1389_l = node1388_l & ~pixel[600];
      node1390_r = node1389_l & pixel[215];
      node1390_l = node1389_l & ~pixel[215];
      node1391_r = node1390_l & pixel[412];
      node1391_l = node1390_l & ~pixel[412];
      node1392 = node1391_l;
      node1393_r = node1391_r & pixel[402];
      node1393_l = node1391_r & ~pixel[402];
      node1394 = node1393_l;
      node1395 = node1393_r;
      node1396_r = node1390_r & pixel[439];
      node1396_l = node1390_r & ~pixel[439];
      node1397_r = node1396_l & pixel[400];
      node1397_l = node1396_l & ~pixel[400];
      node1398 = node1397_l;
      node1399 = node1397_r;
      node1400_r = node1396_r & pixel[208];
      node1400_l = node1396_r & ~pixel[208];
      node1401 = node1400_l;
      node1402 = node1400_r;
      node1403_r = node1389_r & pixel[463];
      node1403_l = node1389_r & ~pixel[463];
      node1404 = node1403_l;
      node1405_r = node1403_r & pixel[689];
      node1405_l = node1403_r & ~pixel[689];
      node1406_r = node1405_l & pixel[455];
      node1406_l = node1405_l & ~pixel[455];
      node1407 = node1406_l;
      node1408 = node1406_r;
      node1409 = node1405_r;
      node1410_r = node1388_r & pixel[371];
      node1410_l = node1388_r & ~pixel[371];
      node1411_r = node1410_l & pixel[204];
      node1411_l = node1410_l & ~pixel[204];
      node1412_r = node1411_l & pixel[577];
      node1412_l = node1411_l & ~pixel[577];
      node1413_r = node1412_l & pixel[566];
      node1413_l = node1412_l & ~pixel[566];
      node1414 = node1413_l;
      node1415 = node1413_r;
      node1416_r = node1412_r & pixel[570];
      node1416_l = node1412_r & ~pixel[570];
      node1417 = node1416_l;
      node1418 = node1416_r;
      node1419_r = node1411_r & pixel[519];
      node1419_l = node1411_r & ~pixel[519];
      node1420_r = node1419_l & pixel[571];
      node1420_l = node1419_l & ~pixel[571];
      node1421 = node1420_l;
      node1422 = node1420_r;
      node1423_r = node1419_r & pixel[604];
      node1423_l = node1419_r & ~pixel[604];
      node1424 = node1423_l;
      node1425 = node1423_r;
      node1426_r = node1410_r & pixel[154];
      node1426_l = node1410_r & ~pixel[154];
      node1427_r = node1426_l & pixel[662];
      node1427_l = node1426_l & ~pixel[662];
      node1428_r = node1427_l & pixel[455];
      node1428_l = node1427_l & ~pixel[455];
      node1429 = node1428_l;
      node1430 = node1428_r;
      node1431 = node1427_r;
      node1432_r = node1426_r & pixel[542];
      node1432_l = node1426_r & ~pixel[542];
      node1433_r = node1432_l & pixel[240];
      node1433_l = node1432_l & ~pixel[240];
      node1434 = node1433_l;
      node1435 = node1433_r;
      node1436 = node1432_r;
      node1437_r = node1387_r & pixel[466];
      node1437_l = node1387_r & ~pixel[466];
      node1438_r = node1437_l & pixel[432];
      node1438_l = node1437_l & ~pixel[432];
      node1439_r = node1438_l & pixel[405];
      node1439_l = node1438_l & ~pixel[405];
      node1440_r = node1439_l & pixel[634];
      node1440_l = node1439_l & ~pixel[634];
      node1441_r = node1440_l & pixel[597];
      node1441_l = node1440_l & ~pixel[597];
      node1442 = node1441_l;
      node1443 = node1441_r;
      node1444_r = node1440_r & pixel[469];
      node1444_l = node1440_r & ~pixel[469];
      node1445 = node1444_l;
      node1446 = node1444_r;
      node1447_r = node1439_r & pixel[524];
      node1447_l = node1439_r & ~pixel[524];
      node1448_r = node1447_l & pixel[606];
      node1448_l = node1447_l & ~pixel[606];
      node1449 = node1448_l;
      node1450 = node1448_r;
      node1451_r = node1447_r & pixel[463];
      node1451_l = node1447_r & ~pixel[463];
      node1452 = node1451_l;
      node1453 = node1451_r;
      node1454_r = node1438_r & pixel[176];
      node1454_l = node1438_r & ~pixel[176];
      node1455_r = node1454_l & pixel[263];
      node1455_l = node1454_l & ~pixel[263];
      node1456_r = node1455_l & pixel[269];
      node1456_l = node1455_l & ~pixel[269];
      node1457 = node1456_l;
      node1458 = node1456_r;
      node1459_r = node1455_r & pixel[636];
      node1459_l = node1455_r & ~pixel[636];
      node1460 = node1459_l;
      node1461 = node1459_r;
      node1462_r = node1454_r & pixel[412];
      node1462_l = node1454_r & ~pixel[412];
      node1463_r = node1462_l & pixel[345];
      node1463_l = node1462_l & ~pixel[345];
      node1464 = node1463_l;
      node1465 = node1463_r;
      node1466_r = node1462_r & pixel[603];
      node1466_l = node1462_r & ~pixel[603];
      node1467 = node1466_l;
      node1468 = node1466_r;
      node1469_r = node1437_r & pixel[489];
      node1469_l = node1437_r & ~pixel[489];
      node1470_r = node1469_l & pixel[546];
      node1470_l = node1469_l & ~pixel[546];
      node1471_r = node1470_l & pixel[431];
      node1471_l = node1470_l & ~pixel[431];
      node1472_r = node1471_l & pixel[377];
      node1472_l = node1471_l & ~pixel[377];
      node1473 = node1472_l;
      node1474 = node1472_r;
      node1475_r = node1471_r & pixel[440];
      node1475_l = node1471_r & ~pixel[440];
      node1476 = node1475_l;
      node1477 = node1475_r;
      node1478_r = node1470_r & pixel[402];
      node1478_l = node1470_r & ~pixel[402];
      node1479_r = node1478_l & pixel[220];
      node1479_l = node1478_l & ~pixel[220];
      node1480 = node1479_l;
      node1481 = node1479_r;
      node1482_r = node1478_r & pixel[572];
      node1482_l = node1478_r & ~pixel[572];
      node1483 = node1482_l;
      node1484 = node1482_r;
      node1485_r = node1469_r & pixel[433];
      node1485_l = node1469_r & ~pixel[433];
      node1486_r = node1485_l & pixel[399];
      node1486_l = node1485_l & ~pixel[399];
      node1487_r = node1486_l & pixel[401];
      node1487_l = node1486_l & ~pixel[401];
      node1488 = node1487_l;
      node1489 = node1487_r;
      node1490_r = node1486_r & pixel[185];
      node1490_l = node1486_r & ~pixel[185];
      node1491 = node1490_l;
      node1492 = node1490_r;
      node1493_r = node1485_r & pixel[155];
      node1493_l = node1485_r & ~pixel[155];
      node1494_r = node1493_l & pixel[454];
      node1494_l = node1493_l & ~pixel[454];
      node1495 = node1494_l;
      node1496 = node1494_r;
      node1497_r = node1493_r & pixel[444];
      node1497_l = node1493_r & ~pixel[444];
      node1498 = node1497_l;
      node1499 = node1497_r;
      node1500_r = node1274_r & pixel[215];
      node1500_l = node1274_r & ~pixel[215];
      node1501_r = node1500_l & pixel[217];
      node1501_l = node1500_l & ~pixel[217];
      node1502_r = node1501_l & pixel[625];
      node1502_l = node1501_l & ~pixel[625];
      node1503_r = node1502_l & pixel[352];
      node1503_l = node1502_l & ~pixel[352];
      node1504_r = node1503_l & pixel[299];
      node1504_l = node1503_l & ~pixel[299];
      node1505_r = node1504_l & pixel[230];
      node1505_l = node1504_l & ~pixel[230];
      node1506_r = node1505_l & pixel[487];
      node1506_l = node1505_l & ~pixel[487];
      node1507 = node1506_l;
      node1508 = node1506_r;
      node1509 = node1505_r;
      node1510_r = node1504_r & pixel[627];
      node1510_l = node1504_r & ~pixel[627];
      node1511 = node1510_l;
      node1512 = node1510_r;
      node1513_r = node1503_r & pixel[297];
      node1513_l = node1503_r & ~pixel[297];
      node1514_r = node1513_l & pixel[508];
      node1514_l = node1513_l & ~pixel[508];
      node1515_r = node1514_l & pixel[150];
      node1515_l = node1514_l & ~pixel[150];
      node1516 = node1515_l;
      node1517 = node1515_r;
      node1518 = node1514_r;
      node1519_r = node1513_r & pixel[264];
      node1519_l = node1513_r & ~pixel[264];
      node1520_r = node1519_l & pixel[289];
      node1520_l = node1519_l & ~pixel[289];
      node1521 = node1520_l;
      node1522 = node1520_r;
      node1523_r = node1519_r & pixel[543];
      node1523_l = node1519_r & ~pixel[543];
      node1524 = node1523_l;
      node1525 = node1523_r;
      node1526_r = node1502_r & pixel[456];
      node1526_l = node1502_r & ~pixel[456];
      node1527_r = node1526_l & pixel[262];
      node1527_l = node1526_l & ~pixel[262];
      node1528_r = node1527_l & pixel[324];
      node1528_l = node1527_l & ~pixel[324];
      node1529_r = node1528_l & pixel[240];
      node1529_l = node1528_l & ~pixel[240];
      node1530 = node1529_l;
      node1531 = node1529_r;
      node1532_r = node1528_r & pixel[485];
      node1532_l = node1528_r & ~pixel[485];
      node1533 = node1532_l;
      node1534 = node1532_r;
      node1535_r = node1527_r & pixel[553];
      node1535_l = node1527_r & ~pixel[553];
      node1536_r = node1535_l & pixel[384];
      node1536_l = node1535_l & ~pixel[384];
      node1537 = node1536_l;
      node1538 = node1536_r;
      node1539 = node1535_r;
      node1540_r = node1526_r & pixel[410];
      node1540_l = node1526_r & ~pixel[410];
      node1541_r = node1540_l & pixel[328];
      node1541_l = node1540_l & ~pixel[328];
      node1542_r = node1541_l & pixel[269];
      node1542_l = node1541_l & ~pixel[269];
      node1543 = node1542_l;
      node1544 = node1542_r;
      node1545 = node1541_r;
      node1546_r = node1540_r & pixel[259];
      node1546_l = node1540_r & ~pixel[259];
      node1547_r = node1546_l & pixel[461];
      node1547_l = node1546_l & ~pixel[461];
      node1548 = node1547_l;
      node1549 = node1547_r;
      node1550_r = node1546_r & pixel[357];
      node1550_l = node1546_r & ~pixel[357];
      node1551 = node1550_l;
      node1552 = node1550_r;
      node1553_r = node1501_r & pixel[621];
      node1553_l = node1501_r & ~pixel[621];
      node1554_r = node1553_l & pixel[602];
      node1554_l = node1553_l & ~pixel[602];
      node1555 = node1554_l;
      node1556_r = node1554_r & pixel[632];
      node1556_l = node1554_r & ~pixel[632];
      node1557_r = node1556_l & pixel[426];
      node1557_l = node1556_l & ~pixel[426];
      node1558 = node1557_l;
      node1559_r = node1557_r & pixel[571];
      node1559_l = node1557_r & ~pixel[571];
      node1560 = node1559_l;
      node1561 = node1559_r;
      node1562 = node1556_r;
      node1563_r = node1553_r & pixel[489];
      node1563_l = node1553_r & ~pixel[489];
      node1564 = node1563_l;
      node1565 = node1563_r;
      node1566_r = node1500_r & pixel[627];
      node1566_l = node1500_r & ~pixel[627];
      node1567_r = node1566_l & pixel[319];
      node1567_l = node1566_l & ~pixel[319];
      node1568_r = node1567_l & pixel[569];
      node1568_l = node1567_l & ~pixel[569];
      node1569_r = node1568_l & pixel[491];
      node1569_l = node1568_l & ~pixel[491];
      node1570 = node1569_l;
      node1571 = node1569_r;
      node1572_r = node1568_r & pixel[412];
      node1572_l = node1568_r & ~pixel[412];
      node1573 = node1572_l;
      node1574_r = node1572_r & pixel[294];
      node1574_l = node1572_r & ~pixel[294];
      node1575 = node1574_l;
      node1576_r = node1574_r & pixel[378];
      node1576_l = node1574_r & ~pixel[378];
      node1577 = node1576_l;
      node1578 = node1576_r;
      node1579_r = node1567_r & pixel[490];
      node1579_l = node1567_r & ~pixel[490];
      node1580_r = node1579_l & pixel[289];
      node1580_l = node1579_l & ~pixel[289];
      node1581 = node1580_l;
      node1582 = node1580_r;
      node1583_r = node1579_r & pixel[629];
      node1583_l = node1579_r & ~pixel[629];
      node1584_r = node1583_l & pixel[247];
      node1584_l = node1583_l & ~pixel[247];
      node1585_r = node1584_l & pixel[624];
      node1585_l = node1584_l & ~pixel[624];
      node1586 = node1585_l;
      node1587 = node1585_r;
      node1588 = node1584_r;
      node1589_r = node1583_r & pixel[297];
      node1589_l = node1583_r & ~pixel[297];
      node1590 = node1589_l;
      node1591 = node1589_r;
      node1592_r = node1566_r & pixel[346];
      node1592_l = node1566_r & ~pixel[346];
      node1593_r = node1592_l & pixel[269];
      node1593_l = node1592_l & ~pixel[269];
      node1594_r = node1593_l & pixel[375];
      node1594_l = node1593_l & ~pixel[375];
      node1595_r = node1594_l & pixel[274];
      node1595_l = node1594_l & ~pixel[274];
      node1596 = node1595_l;
      node1597_r = node1595_r & pixel[464];
      node1597_l = node1595_r & ~pixel[464];
      node1598 = node1597_l;
      node1599 = node1597_r;
      node1600_r = node1594_r & pixel[541];
      node1600_l = node1594_r & ~pixel[541];
      node1601 = node1600_l;
      node1602 = node1600_r;
      node1603_r = node1593_r & pixel[320];
      node1603_l = node1593_r & ~pixel[320];
      node1604_r = node1603_l & pixel[453];
      node1604_l = node1603_l & ~pixel[453];
      node1605_r = node1604_l & pixel[635];
      node1605_l = node1604_l & ~pixel[635];
      node1606 = node1605_l;
      node1607 = node1605_r;
      node1608_r = node1604_r & pixel[620];
      node1608_l = node1604_r & ~pixel[620];
      node1609 = node1608_l;
      node1610 = node1608_r;
      node1611_r = node1603_r & pixel[628];
      node1611_l = node1603_r & ~pixel[628];
      node1612 = node1611_l;
      node1613_r = node1611_r & pixel[127];
      node1613_l = node1611_r & ~pixel[127];
      node1614 = node1613_l;
      node1615 = node1613_r;
      node1616_r = node1592_r & pixel[327];
      node1616_l = node1592_r & ~pixel[327];
      node1617_r = node1616_l & pixel[235];
      node1617_l = node1616_l & ~pixel[235];
      node1618_r = node1617_l & pixel[270];
      node1618_l = node1617_l & ~pixel[270];
      node1619 = node1618_l;
      node1620 = node1618_r;
      node1621 = node1617_r;
      node1622_r = node1616_r & pixel[406];
      node1622_l = node1616_r & ~pixel[406];
      node1623_r = node1622_l & pixel[236];
      node1623_l = node1622_l & ~pixel[236];
      node1624 = node1623_l;
      node1625_r = node1623_r & pixel[609];
      node1625_l = node1623_r & ~pixel[609];
      node1626 = node1625_l;
      node1627 = node1625_r;
      node1628_r = node1622_r & pixel[317];
      node1628_l = node1622_r & ~pixel[317];
      node1629_r = node1628_l & pixel[428];
      node1629_l = node1628_l & ~pixel[428];
      node1630 = node1629_l;
      node1631 = node1629_r;
      node1632 = node1628_r;
      result0 = node13 | node18 | node21 | node29 | node41 | node47 | node55 | node57 | node61 | node67 | node77 | node82 | node83 | node91 | node96 | node99 | node100 | node103 | node107 | node118 | node119 | node131 | node137 | node142 | node149 | node150 | node152 | node157 | node161 | node165 | node167 | node174 | node175 | node177 | node183 | node184 | node187 | node193 | node194 | node201 | node297 | node313 | node346 | node372 | node374 | node398 | node411 | node500 | node503 | node607 | node609 | node653 | node654 | node657 | node681 | node686 | node776 | node809 | node1045 | node1048 | node1089 | node1103 | node1104 | node1129 | node1136 | node1147 | node1154 | node1155 | node1237 | node1300 | node1331 | node1353 | node1382 | node1446 | node1473 | node1483 | node1484 | node1524 | node1561 | node1588 | node1626 | node1631;
      result1 = node225 | node232 | node421 | node425 | node431 | node439 | node444 | node452 | node453 | node459 | node467 | node471 | node474 | node622 | node628 | node663 | node722 | node725 | node729 | node879 | node1184 | node1249 | node1262 | node1289 | node1533;
      result2 = node14 | node33 | node42 | node54 | node68 | node78 | node86 | node104 | node120 | node168 | node213 | node216 | node242 | node243 | node247 | node248 | node250 | node264 | node272 | node273 | node277 | node278 | node281 | node293 | node305 | node379 | node397 | node402 | node422 | node477 | node554 | node577 | node578 | node580 | node587 | node634 | node694 | node695 | node698 | node712 | node714 | node732 | node743 | node747 | node752 | node755 | node760 | node763 | node773 | node782 | node789 | node801 | node802 | node812 | node815 | node833 | node843 | node850 | node895 | node909 | node926 | node970 | node978 | node994 | node995 | node999 | node1001 | node1059 | node1064 | node1070 | node1113 | node1116 | node1128 | node1131 | node1132 | node1138 | node1145 | node1151 | node1166 | node1169 | node1178 | node1252 | node1257 | node1270 | node1272 | node1282 | node1283 | node1286 | node1290 | node1293 | node1324 | node1345 | node1346 | node1354 | node1358 | node1367 | node1371 | node1376 | node1385 | node1445 | node1453 | node1464 | node1499 | node1512 | node1521 | node1534 | node1544 | node1555 | node1560 | node1565 | node1571 | node1573 | node1575 | node1578 | node1586 | node1587 | node1596 | node1599 | node1602 | node1606 | node1607 | node1610 | node1612 | node1627;
      result3 = node17 | node20 | node58 | node60 | node70 | node89 | node90 | node228 | node283 | node321 | node324 | node368 | node369 | node401 | node470 | node526 | node546 | node549 | node562 | node568 | node569 | node571 | node604 | node629 | node640 | node648 | node651 | node664 | node666 | node670 | node673 | node674 | node678 | node682 | node688 | node708 | node709 | node721 | node737 | node739 | node740 | node783 | node786 | node797 | node825 | node836 | node848 | node856 | node857 | node863 | node864 | node866 | node894 | node967 | node977 | node1006 | node1009 | node1014 | node1030 | node1033 | node1060 | node1063 | node1069 | node1074 | node1075 | node1078 | node1084 | node1091 | node1114 | node1152 | node1193 | node1195 | node1196 | node1198 | node1202 | node1204 | node1207 | node1210 | node1219 | node1221 | node1222 | node1225 | node1226 | node1229 | node1236 | node1240 | node1241 | node1244 | node1266 | node1269 | node1273 | node1373 | node1378 | node1386 | node1417 | node1421 | node1425 | node1435 | node1452 | node1474 | node1564 | node1577 | node1581 | node1598 | node1609 | node1615 | node1620 | node1630;
      result4 = node112 | node220 | node254 | node267 | node290 | node292 | node296 | node299 | node337 | node345 | node353 | node358 | node378 | node394 | node406 | node412 | node440 | node484 | node531 | node547 | node553 | node556 | node596 | node605 | node901 | node916 | node917 | node924 | node934 | node937 | node941 | node944 | node949 | node950 | node952 | node953 | node956 | node972 | node976 | node982 | node984 | node1016 | node1025 | node1029 | node1038 | node1044 | node1071 | node1077 | node1099 | node1139 | node1177 | node1180 | node1181 | node1185 | node1297 | node1301 | node1316 | node1320 | node1321 | node1328 | node1335 | node1395 | node1401 | node1407 | node1408 | node1481 | node1491 | node1496 | node1522 | node1582 | node1591;
      result5 = node11 | node26 | node32 | node35 | node44 | node45 | node50 | node71 | node75 | node97 | node106 | node115 | node127 | node135 | node143 | node145 | node164 | node191 | node199 | node210 | node212 | node217 | node219 | node227 | node231 | node279 | node284 | node289 | node306 | node309 | node312 | node320 | node331 | node332 | node343 | node351 | node356 | node365 | node373 | node381 | node385 | node388 | node389 | node436 | node446 | node455 | node462 | node491 | node499 | node506 | node509 | node518 | node522 | node535 | node585 | node621 | node625 | node626 | node633 | node637 | node647 | node667 | node671 | node679 | node685 | node689 | node706 | node713 | node736 | node798 | node806 | node814 | node826 | node829 | node835 | node859 | node867 | node888 | node892 | node923 | node927 | node942 | node965 | node966 | node985 | node998 | node1013 | node1017 | node1037 | node1040 | node1041 | node1047 | node1056 | node1083 | node1086 | node1087 | node1096 | node1107 | node1160 | node1163 | node1188 | node1192 | node1212 | node1218 | node1228 | node1233 | node1234 | node1243 | node1263 | node1379 | node1392 | node1399 | node1434 | node1518 | node1539 | node1551 | node1558;
      result6 = node25 | node28 | node74 | node111 | node128 | node138 | node146 | node186 | node190 | node209 | node233 | node238 | node239 | node265 | node271 | node310 | node327 | node338 | node340 | node350 | node354 | node359 | node366 | node386 | node409 | node478 | node494 | node495 | node525 | node532 | node561 | node564 | node588 | node595 | node598 | node603 | node636 | node697 | node701 | node731 | node753 | node768 | node769 | node772 | node792 | node807 | node810 | node891 | node896 | node902 | node935 | node1057 | node1106 | node1117 | node1121 | node1135 | node1144 | node1159 | node1162 | node1298 | node1304 | node1307 | node1314 | node1317 | node1347 | node1350 | node1351 | node1357 | node1359 | node1364 | node1365 | node1368 | node1372 | node1383 | node1507 | node1508 | node1511 | node1516 | node1517 | node1525 | node1530 | node1531 | node1538 | node1543 | node1545 | node1548 | node1549 | node1552 | node1562 | node1570 | node1590 | node1601 | node1614 | node1619 | node1621 | node1624 | node1632;
      result7 = node10 | node36 | node49 | node130 | node134 | node156 | node162 | node179 | node197 | node224 | node258 | node428 | node432 | node460 | node485 | node565 | node572 | node581 | node589 | node599 | node618 | node649 | node828 | node832 | node840 | node841 | node847 | node871 | node887 | node905 | node945 | node957 | node960 | node981 | node1258 | node1285 | node1394 | node1424 | node1429 | node1442 | node1488;
      result8 = node114 | node153 | node241 | node251 | node257 | node268 | node300 | node323 | node330 | node341 | node382 | node424 | node429 | node437 | node443 | node456 | node463 | node468 | node475 | node488 | node492 | node502 | node507 | node510 | node515 | node516 | node519 | node523 | node530 | node536 | node538 | node539 | node557 | node641 | node642 | node656 | node705 | node724 | node728 | node744 | node746 | node756 | node759 | node762 | node775 | node785 | node790 | node793 | node800 | node844 | node875 | node878 | node881 | node882 | node971 | node1026 | node1032 | node1065 | node1092 | node1100 | node1123 | node1148 | node1167 | node1170 | node1187 | node1205 | node1211 | node1253 | node1256 | node1265 | node1292 | node1305 | node1308 | node1323 | node1332 | node1398 | node1402 | node1404 | node1409 | node1414 | node1415 | node1418 | node1422 | node1431 | node1436 | node1443 | node1449 | node1450 | node1457 | node1458 | node1460 | node1461 | node1465 | node1467 | node1468 | node1476 | node1477 | node1480 | node1489 | node1495 | node1498 | node1509 | node1537;
      result9 = node85 | node178 | node200 | node255 | node304 | node328 | node395 | node403 | node408 | node447 | node487 | node550 | node584 | node593 | node610 | node619 | node700 | node767 | node851 | node860 | node872 | node874 | node904 | node908 | node911 | node912 | node919 | node920 | node938 | node959 | node991 | node992 | node1002 | node1007 | node1010 | node1022 | node1023 | node1097 | node1120 | node1124 | node1199 | node1250 | node1313 | node1329 | node1336 | node1338 | node1339 | node1430 | node1492;

      tree_9 = {result9, result8, result7, result6, result5, result4, result3, result2, result1, result0};
    end
  endfunction

  wire [9:0] res_tree_0;
  assign res_tree_0 = tree_0(image);
  wire [9:0] res_tree_1;
  assign res_tree_1 = tree_1(image);
  wire [9:0] res_tree_2;
  assign res_tree_2 = tree_2(image);
  wire [9:0] res_tree_3;
  assign res_tree_3 = tree_3(image);
  wire [9:0] res_tree_4;
  assign res_tree_4 = tree_4(image);
  wire [9:0] res_tree_5;
  assign res_tree_5 = tree_5(image);
  wire [9:0] res_tree_6;
  assign res_tree_6 = tree_6(image);
  wire [9:0] res_tree_7;
  assign res_tree_7 = tree_7(image);
  wire [9:0] res_tree_8;
  assign res_tree_8 = tree_8(image);
  wire [9:0] res_tree_9;
  assign res_tree_9 = tree_9(image);

  wire [7:0] res_sum_0;
  assign res_sum_0 = {7'b0000000, res_tree_0[0]} + {7'b0000000, res_tree_1[0]} + {7'b0000000, res_tree_2[0]} + {7'b0000000, res_tree_3[0]} + {7'b0000000, res_tree_4[0]} + {7'b0000000, res_tree_5[0]} + {7'b0000000, res_tree_6[0]} + {7'b0000000, res_tree_7[0]} + {7'b0000000, res_tree_8[0]} + {7'b0000000, res_tree_9[0]};
  wire [7:0] res_sum_1;
  assign res_sum_1 = {7'b0000000, res_tree_0[1]} + {7'b0000000, res_tree_1[1]} + {7'b0000000, res_tree_2[1]} + {7'b0000000, res_tree_3[1]} + {7'b0000000, res_tree_4[1]} + {7'b0000000, res_tree_5[1]} + {7'b0000000, res_tree_6[1]} + {7'b0000000, res_tree_7[1]} + {7'b0000000, res_tree_8[1]} + {7'b0000000, res_tree_9[1]};
  wire [7:0] res_sum_2;
  assign res_sum_2 = {7'b0000000, res_tree_0[2]} + {7'b0000000, res_tree_1[2]} + {7'b0000000, res_tree_2[2]} + {7'b0000000, res_tree_3[2]} + {7'b0000000, res_tree_4[2]} + {7'b0000000, res_tree_5[2]} + {7'b0000000, res_tree_6[2]} + {7'b0000000, res_tree_7[2]} + {7'b0000000, res_tree_8[2]} + {7'b0000000, res_tree_9[2]};
  wire [7:0] res_sum_3;
  assign res_sum_3 = {7'b0000000, res_tree_0[3]} + {7'b0000000, res_tree_1[3]} + {7'b0000000, res_tree_2[3]} + {7'b0000000, res_tree_3[3]} + {7'b0000000, res_tree_4[3]} + {7'b0000000, res_tree_5[3]} + {7'b0000000, res_tree_6[3]} + {7'b0000000, res_tree_7[3]} + {7'b0000000, res_tree_8[3]} + {7'b0000000, res_tree_9[3]};
  wire [7:0] res_sum_4;
  assign res_sum_4 = {7'b0000000, res_tree_0[4]} + {7'b0000000, res_tree_1[4]} + {7'b0000000, res_tree_2[4]} + {7'b0000000, res_tree_3[4]} + {7'b0000000, res_tree_4[4]} + {7'b0000000, res_tree_5[4]} + {7'b0000000, res_tree_6[4]} + {7'b0000000, res_tree_7[4]} + {7'b0000000, res_tree_8[4]} + {7'b0000000, res_tree_9[4]};
  wire [7:0] res_sum_5;
  assign res_sum_5 = {7'b0000000, res_tree_0[5]} + {7'b0000000, res_tree_1[5]} + {7'b0000000, res_tree_2[5]} + {7'b0000000, res_tree_3[5]} + {7'b0000000, res_tree_4[5]} + {7'b0000000, res_tree_5[5]} + {7'b0000000, res_tree_6[5]} + {7'b0000000, res_tree_7[5]} + {7'b0000000, res_tree_8[5]} + {7'b0000000, res_tree_9[5]};
  wire [7:0] res_sum_6;
  assign res_sum_6 = {7'b0000000, res_tree_0[6]} + {7'b0000000, res_tree_1[6]} + {7'b0000000, res_tree_2[6]} + {7'b0000000, res_tree_3[6]} + {7'b0000000, res_tree_4[6]} + {7'b0000000, res_tree_5[6]} + {7'b0000000, res_tree_6[6]} + {7'b0000000, res_tree_7[6]} + {7'b0000000, res_tree_8[6]} + {7'b0000000, res_tree_9[6]};
  wire [7:0] res_sum_7;
  assign res_sum_7 = {7'b0000000, res_tree_0[7]} + {7'b0000000, res_tree_1[7]} + {7'b0000000, res_tree_2[7]} + {7'b0000000, res_tree_3[7]} + {7'b0000000, res_tree_4[7]} + {7'b0000000, res_tree_5[7]} + {7'b0000000, res_tree_6[7]} + {7'b0000000, res_tree_7[7]} + {7'b0000000, res_tree_8[7]} + {7'b0000000, res_tree_9[7]};
  wire [7:0] res_sum_8;
  assign res_sum_8 = {7'b0000000, res_tree_0[8]} + {7'b0000000, res_tree_1[8]} + {7'b0000000, res_tree_2[8]} + {7'b0000000, res_tree_3[8]} + {7'b0000000, res_tree_4[8]} + {7'b0000000, res_tree_5[8]} + {7'b0000000, res_tree_6[8]} + {7'b0000000, res_tree_7[8]} + {7'b0000000, res_tree_8[8]} + {7'b0000000, res_tree_9[8]};
  wire [7:0] res_sum_9;
  assign res_sum_9 = {7'b0000000, res_tree_0[9]} + {7'b0000000, res_tree_1[9]} + {7'b0000000, res_tree_2[9]} + {7'b0000000, res_tree_3[9]} + {7'b0000000, res_tree_4[9]} + {7'b0000000, res_tree_5[9]} + {7'b0000000, res_tree_6[9]} + {7'b0000000, res_tree_7[9]} + {7'b0000000, res_tree_8[9]} + {7'b0000000, res_tree_9[9]};

  wire [7:0] winner_cnt_0vs1;
  wire [7:0] winner_cnt_2vs3;
  wire [7:0] winner_cnt_4vs5;
    wire [7:0] winner_cnt_6vs7;
    wire [7:0] winner_cnt_8vs9;
    wire [7:0] winner_cnt_01vs23;
    wire [7:0] winner_cnt_45vs67;
    wire [7:0] winner_cnt_0123vs4567;

    wire [3:0] winner_0vs1;
    wire [3:0] winner_2vs3;
    wire [3:0] winner_4vs5;
    wire [3:0] winner_6vs7;
    wire [3:0] winner_8vs9;
    wire [3:0] winner_01vs23;
    wire [3:0] winner_45vs67;
    wire [3:0] winner_0123vs4567;
    wire [3:0] winner;

  assign winner_cnt_0vs1 = res_sum_1 > res_sum_0 ? res_sum_1 : res_sum_0;
  assign winner_0vs1     = res_sum_1 > res_sum_0 ? 1 : 0;
  assign winner_cnt_2vs3 = res_sum_3 > res_sum_2 ? res_sum_3 : res_sum_2;
  assign winner_2vs3     = res_sum_3 > res_sum_2 ? 3 : 2;
  assign winner_cnt_4vs5 = res_sum_5 > res_sum_4 ? res_sum_5 : res_sum_4;
  assign winner_4vs5     = res_sum_5 > res_sum_4 ? 5 : 4;
  assign winner_cnt_6vs7 = res_sum_7 > res_sum_6 ? res_sum_7 : res_sum_6;
  assign winner_6vs7     = res_sum_7 > res_sum_6 ? 7 : 6;
  assign winner_cnt_8vs9 = res_sum_9 > res_sum_8 ? res_sum_9 : res_sum_8;
  assign winner_8vs9     = res_sum_9 > res_sum_8 ? 9 : 8;

  assign winner_cnt_01vs23 = winner_cnt_2vs3 > winner_cnt_0vs1 ? winner_cnt_2vs3 : winner_cnt_0vs1;
  assign winner_01vs23     = winner_cnt_2vs3 > winner_cnt_0vs1 ? winner_2vs3 : winner_0vs1;
  assign winner_cnt_45vs67 = winner_cnt_6vs7 > winner_cnt_4vs5 ? winner_cnt_6vs7 : winner_cnt_4vs5;
  assign winner_45vs67     = winner_cnt_6vs7 > winner_cnt_4vs5 ? winner_6vs7 : winner_4vs5;

  assign winner_cnt_0123vs4567 = winner_cnt_45vs67 > winner_cnt_01vs23 ? winner_cnt_45vs67 : winner_cnt_01vs23;
  assign winner_0123vs4567     = winner_cnt_45vs67 > winner_cnt_01vs23 ? winner_45vs67 : winner_01vs23;

  assign winner = winner_cnt_8vs9 > winner_cnt_0123vs4567 ? winner_8vs9 : winner_0123vs4567;
  assign result = winner;

endmodule
